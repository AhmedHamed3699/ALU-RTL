module sequential_multiplier (A,
    B,
    Product);
 input [31:0] A;
 input [31:0] B;
 output [63:0] Product;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;

 sky130_fd_sc_hd__inv_16 _14469_ (.A(net33),
    .Y(_03178_));
 sky130_fd_sc_hd__inv_16 _14470_ (.A(net1),
    .Y(_03289_));
 sky130_fd_sc_hd__clkinv_16 _14471_ (.A(net25),
    .Y(_03399_));
 sky130_fd_sc_hd__inv_4 _14472_ (.A(net23),
    .Y(_03510_));
 sky130_fd_sc_hd__clkinv_8 _14473_ (.A(net26),
    .Y(_03621_));
 sky130_fd_sc_hd__inv_2 _14474_ (.A(net27),
    .Y(_03731_));
 sky130_fd_sc_hd__inv_2 _14475_ (.A(net28),
    .Y(_03841_));
 sky130_fd_sc_hd__clkinv_4 _14476_ (.A(net29),
    .Y(_03952_));
 sky130_fd_sc_hd__inv_2 _14477_ (.A(net30),
    .Y(_04062_));
 sky130_fd_sc_hd__inv_2 _14478_ (.A(net32),
    .Y(_04172_));
 sky130_fd_sc_hd__inv_2 _14479_ (.A(net2),
    .Y(_04282_));
 sky130_fd_sc_hd__clkinv_4 _14480_ (.A(net3),
    .Y(_04392_));
 sky130_fd_sc_hd__inv_2 _14481_ (.A(net4),
    .Y(_04503_));
 sky130_fd_sc_hd__nand2_1 _14482_ (.A(net33),
    .B(net1),
    .Y(_04613_));
 sky130_fd_sc_hd__inv_2 _14483_ (.A(_04613_),
    .Y(net65));
 sky130_fd_sc_hd__nor2_8 _14484_ (.A(net409),
    .B(_03399_),
    .Y(_04832_));
 sky130_fd_sc_hd__and2_4 _14485_ (.A(_03399_),
    .B(net409),
    .X(_04942_));
 sky130_fd_sc_hd__nor2_8 _14486_ (.A(_04832_),
    .B(_04942_),
    .Y(_05051_));
 sky130_fd_sc_hd__or2_4 _14487_ (.A(_04832_),
    .B(_04942_),
    .X(_05119_));
 sky130_fd_sc_hd__a21oi_4 _14488_ (.A1(net33),
    .A2(net409),
    .B1(net44),
    .Y(_05130_));
 sky130_fd_sc_hd__a21o_4 _14489_ (.A1(net33),
    .A2(net409),
    .B1(net44),
    .X(_05141_));
 sky130_fd_sc_hd__and3_4 _14490_ (.A(net33),
    .B(net44),
    .C(net409),
    .X(_05152_));
 sky130_fd_sc_hd__nand3_4 _14491_ (.A(net33),
    .B(net44),
    .C(net409),
    .Y(_05163_));
 sky130_fd_sc_hd__nor2_8 _14492_ (.A(net408),
    .B(_05152_),
    .Y(_05174_));
 sky130_fd_sc_hd__nand2_8 _14493_ (.A(_05141_),
    .B(_05163_),
    .Y(_05185_));
 sky130_fd_sc_hd__a21oi_4 _14494_ (.A1(net1),
    .A2(net25),
    .B1(net12),
    .Y(_05196_));
 sky130_fd_sc_hd__a21o_4 _14495_ (.A1(net1),
    .A2(net25),
    .B1(net12),
    .X(_05207_));
 sky130_fd_sc_hd__and3_4 _14496_ (.A(net12),
    .B(net1),
    .C(net25),
    .X(_05218_));
 sky130_fd_sc_hd__nand3_4 _14497_ (.A(net12),
    .B(net1),
    .C(net25),
    .Y(_05229_));
 sky130_fd_sc_hd__nor2_8 _14498_ (.A(net407),
    .B(_05218_),
    .Y(_05239_));
 sky130_fd_sc_hd__nand2_8 _14499_ (.A(_05207_),
    .B(_05229_),
    .Y(_05250_));
 sky130_fd_sc_hd__and3_1 _14500_ (.A(_05207_),
    .B(_05229_),
    .C(net33),
    .X(_05261_));
 sky130_fd_sc_hd__a31o_1 _14501_ (.A1(net1),
    .A2(_05141_),
    .A3(_05163_),
    .B1(_05261_),
    .X(_05272_));
 sky130_fd_sc_hd__or4_1 _14502_ (.A(net408),
    .B(_05152_),
    .C(_05196_),
    .D(_05218_),
    .X(_05283_));
 sky130_fd_sc_hd__o21ai_1 _14503_ (.A1(_04613_),
    .A2(_05283_),
    .B1(_05272_),
    .Y(_05294_));
 sky130_fd_sc_hd__o31a_1 _14504_ (.A1(_03178_),
    .A2(_03289_),
    .A3(_05051_),
    .B1(_05294_),
    .X(_05305_));
 sky130_fd_sc_hd__a41oi_1 _14505_ (.A1(net65),
    .A2(_05119_),
    .A3(_05272_),
    .A4(_05283_),
    .B1(_05305_),
    .Y(net76));
 sky130_fd_sc_hd__o22a_1 _14506_ (.A1(_04832_),
    .A2(_04942_),
    .B1(net65),
    .B2(_05272_),
    .X(_05326_));
 sky130_fd_sc_hd__or2_4 _14507_ (.A(net33),
    .B(net44),
    .X(_05337_));
 sky130_fd_sc_hd__and3b_4 _14508_ (.A_N(net55),
    .B(_05337_),
    .C(net409),
    .X(_05348_));
 sky130_fd_sc_hd__nand3b_4 _14509_ (.A_N(net55),
    .B(_05337_),
    .C(net409),
    .Y(_05359_));
 sky130_fd_sc_hd__a21boi_4 _14510_ (.A1(_05337_),
    .A2(net409),
    .B1_N(net55),
    .Y(_05370_));
 sky130_fd_sc_hd__a21bo_4 _14511_ (.A1(_05337_),
    .A2(net409),
    .B1_N(net55),
    .X(_05381_));
 sky130_fd_sc_hd__nor2_8 _14512_ (.A(net402),
    .B(net399),
    .Y(_05392_));
 sky130_fd_sc_hd__nand2_8 _14513_ (.A(_05359_),
    .B(_05381_),
    .Y(_05403_));
 sky130_fd_sc_hd__nor2_8 _14514_ (.A(net12),
    .B(net1),
    .Y(_05414_));
 sky130_fd_sc_hd__or2_1 _14515_ (.A(net12),
    .B(net1),
    .X(_05425_));
 sky130_fd_sc_hd__o21ai_1 _14516_ (.A1(net12),
    .A2(net1),
    .B1(net25),
    .Y(_05436_));
 sky130_fd_sc_hd__and3_4 _14517_ (.A(_05425_),
    .B(net25),
    .C(_03510_),
    .X(_05447_));
 sky130_fd_sc_hd__o211ai_4 _14518_ (.A1(net12),
    .A2(net1),
    .B1(net25),
    .C1(_03510_),
    .Y(_05458_));
 sky130_fd_sc_hd__o21a_4 _14519_ (.A1(_03399_),
    .A2(_05414_),
    .B1(net23),
    .X(_05469_));
 sky130_fd_sc_hd__nand2_4 _14520_ (.A(_05436_),
    .B(net23),
    .Y(_05480_));
 sky130_fd_sc_hd__o21ai_4 _14521_ (.A1(net12),
    .A2(net1),
    .B1(net23),
    .Y(_05491_));
 sky130_fd_sc_hd__o211a_4 _14522_ (.A1(net12),
    .A2(net1),
    .B1(net25),
    .C1(net23),
    .X(_05501_));
 sky130_fd_sc_hd__or3_4 _14523_ (.A(_03399_),
    .B(_03510_),
    .C(_05414_),
    .X(_05512_));
 sky130_fd_sc_hd__o21a_4 _14524_ (.A1(_03399_),
    .A2(_05414_),
    .B1(_03510_),
    .X(_05523_));
 sky130_fd_sc_hd__o21ai_4 _14525_ (.A1(_03399_),
    .A2(_05414_),
    .B1(_03510_),
    .Y(_05534_));
 sky130_fd_sc_hd__o21ai_4 _14526_ (.A1(_03399_),
    .A2(_05491_),
    .B1(net396),
    .Y(_05545_));
 sky130_fd_sc_hd__nand2_8 _14527_ (.A(_05458_),
    .B(_05480_),
    .Y(_05556_));
 sky130_fd_sc_hd__o211ai_4 _14528_ (.A1(_03399_),
    .A2(_05491_),
    .B1(net33),
    .C1(_05534_),
    .Y(_05567_));
 sky130_fd_sc_hd__a32o_1 _14529_ (.A1(net404),
    .A2(net403),
    .A3(_04613_),
    .B1(_05556_),
    .B2(net33),
    .X(_05578_));
 sky130_fd_sc_hd__or4_1 _14530_ (.A(net65),
    .B(_05185_),
    .C(_05250_),
    .D(_05567_),
    .X(_05589_));
 sky130_fd_sc_hd__o2bb2a_1 _14531_ (.A1_N(_05578_),
    .A2_N(_05589_),
    .B1(_03289_),
    .B2(_05392_),
    .X(_05600_));
 sky130_fd_sc_hd__a31o_1 _14532_ (.A1(net1),
    .A2(net388),
    .A3(_05578_),
    .B1(_05600_),
    .X(_05611_));
 sky130_fd_sc_hd__xnor2_1 _14533_ (.A(_05326_),
    .B(_05611_),
    .Y(net87));
 sky130_fd_sc_hd__a31o_1 _14534_ (.A1(_04613_),
    .A2(_05611_),
    .A3(_05294_),
    .B1(_05051_),
    .X(_05632_));
 sky130_fd_sc_hd__o21ai_4 _14535_ (.A1(net55),
    .A2(_05337_),
    .B1(net409),
    .Y(_05643_));
 sky130_fd_sc_hd__o311a_4 _14536_ (.A1(net33),
    .A2(net44),
    .A3(net55),
    .B1(net58),
    .C1(net409),
    .X(_05654_));
 sky130_fd_sc_hd__and2b_4 _14537_ (.A_N(net58),
    .B(_05643_),
    .X(_05665_));
 sky130_fd_sc_hd__nor2_8 _14538_ (.A(net58),
    .B(_05643_),
    .Y(_05676_));
 sky130_fd_sc_hd__or2_4 _14539_ (.A(net58),
    .B(_05643_),
    .X(_05687_));
 sky130_fd_sc_hd__and2_4 _14540_ (.A(_05643_),
    .B(net58),
    .X(_05698_));
 sky130_fd_sc_hd__nand2_8 _14541_ (.A(_05643_),
    .B(net58),
    .Y(_05709_));
 sky130_fd_sc_hd__nor2_8 _14542_ (.A(_05654_),
    .B(_05665_),
    .Y(_05720_));
 sky130_fd_sc_hd__nor2_8 _14543_ (.A(net384),
    .B(net383),
    .Y(_05731_));
 sky130_fd_sc_hd__nand2_2 _14544_ (.A(_05578_),
    .B(net1),
    .Y(_05742_));
 sky130_fd_sc_hd__nor3_4 _14545_ (.A(net12),
    .B(net1),
    .C(net23),
    .Y(_05753_));
 sky130_fd_sc_hd__o311a_4 _14546_ (.A1(net12),
    .A2(net1),
    .A3(net23),
    .B1(_03621_),
    .C1(net25),
    .X(_05763_));
 sky130_fd_sc_hd__o311ai_4 _14547_ (.A1(net12),
    .A2(net1),
    .A3(net23),
    .B1(_03621_),
    .C1(net25),
    .Y(_05774_));
 sky130_fd_sc_hd__o21a_4 _14548_ (.A1(_03399_),
    .A2(_05753_),
    .B1(net26),
    .X(_05785_));
 sky130_fd_sc_hd__o21ai_4 _14549_ (.A1(_03399_),
    .A2(_05753_),
    .B1(net26),
    .Y(_05796_));
 sky130_fd_sc_hd__o311a_4 _14550_ (.A1(net12),
    .A2(net1),
    .A3(net23),
    .B1(net26),
    .C1(net25),
    .X(_05807_));
 sky130_fd_sc_hd__o311ai_4 _14551_ (.A1(net12),
    .A2(net1),
    .A3(net23),
    .B1(net26),
    .C1(net25),
    .Y(_05818_));
 sky130_fd_sc_hd__o21a_4 _14552_ (.A1(_03399_),
    .A2(_05753_),
    .B1(_03621_),
    .X(_05829_));
 sky130_fd_sc_hd__o21bai_4 _14553_ (.A1(_03399_),
    .A2(_05753_),
    .B1_N(net26),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_8 _14554_ (.A(net406),
    .B(_05840_),
    .Y(_05851_));
 sky130_fd_sc_hd__nand2_8 _14555_ (.A(net395),
    .B(_05796_),
    .Y(_05862_));
 sky130_fd_sc_hd__nand3_2 _14556_ (.A(_05840_),
    .B(net33),
    .C(_05818_),
    .Y(_05873_));
 sky130_fd_sc_hd__a31oi_2 _14557_ (.A1(_05840_),
    .A2(net33),
    .A3(_05818_),
    .B1(_05556_),
    .Y(_05884_));
 sky130_fd_sc_hd__o21ai_4 _14558_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_05873_),
    .Y(_05895_));
 sky130_fd_sc_hd__a41oi_2 _14559_ (.A1(_05556_),
    .A2(_05818_),
    .A3(_05840_),
    .A4(net33),
    .B1(_05185_),
    .Y(_05906_));
 sky130_fd_sc_hd__a41o_1 _14560_ (.A1(_05556_),
    .A2(_05818_),
    .A3(_05840_),
    .A4(net33),
    .B1(_05185_),
    .X(_05917_));
 sky130_fd_sc_hd__nand2_1 _14561_ (.A(_05906_),
    .B(_05895_),
    .Y(_05928_));
 sky130_fd_sc_hd__o2111ai_2 _14562_ (.A1(net408),
    .A2(_05152_),
    .B1(net33),
    .C1(_05818_),
    .D1(_05840_),
    .Y(_05939_));
 sky130_fd_sc_hd__nand3_2 _14563_ (.A(_03289_),
    .B(_05458_),
    .C(_05480_),
    .Y(_05950_));
 sky130_fd_sc_hd__nand2_2 _14564_ (.A(_05950_),
    .B(_05261_),
    .Y(_05961_));
 sky130_fd_sc_hd__nand4_1 _14565_ (.A(_05950_),
    .B(net403),
    .C(net404),
    .D(net33),
    .Y(_05972_));
 sky130_fd_sc_hd__a22oi_2 _14566_ (.A1(_05939_),
    .A2(_05972_),
    .B1(_05906_),
    .B2(_05895_),
    .Y(_05983_));
 sky130_fd_sc_hd__o2bb2ai_1 _14567_ (.A1_N(_05939_),
    .A2_N(_05972_),
    .B1(_05884_),
    .B2(_05917_),
    .Y(_05994_));
 sky130_fd_sc_hd__o2111a_1 _14568_ (.A1(_05567_),
    .A2(_05851_),
    .B1(_05961_),
    .C1(net404),
    .D1(_05895_),
    .X(_06004_));
 sky130_fd_sc_hd__o2111ai_4 _14569_ (.A1(_05567_),
    .A2(_05851_),
    .B1(_05961_),
    .C1(net404),
    .D1(_05895_),
    .Y(_06015_));
 sky130_fd_sc_hd__nand2_2 _14570_ (.A(_05994_),
    .B(_06015_),
    .Y(_06026_));
 sky130_fd_sc_hd__a21oi_2 _14571_ (.A1(_05994_),
    .A2(_06015_),
    .B1(_05250_),
    .Y(_06037_));
 sky130_fd_sc_hd__o21bai_4 _14572_ (.A1(_05983_),
    .A2(_06004_),
    .B1_N(_05250_),
    .Y(_06048_));
 sky130_fd_sc_hd__o22a_1 _14573_ (.A1(_05196_),
    .A2(_05218_),
    .B1(net404),
    .B2(_05873_),
    .X(_06059_));
 sky130_fd_sc_hd__a21oi_1 _14574_ (.A1(_05928_),
    .A2(_06059_),
    .B1(_06037_),
    .Y(_06070_));
 sky130_fd_sc_hd__a22o_1 _14575_ (.A1(_05928_),
    .A2(_06059_),
    .B1(_06026_),
    .B2(net403),
    .X(_06081_));
 sky130_fd_sc_hd__o211ai_4 _14576_ (.A1(net402),
    .A2(net399),
    .B1(_05742_),
    .C1(_06081_),
    .Y(_06092_));
 sky130_fd_sc_hd__nand4_2 _14577_ (.A(net388),
    .B(_06070_),
    .C(_05578_),
    .D(net1),
    .Y(_06103_));
 sky130_fd_sc_hd__a21oi_2 _14578_ (.A1(_05928_),
    .A2(_06059_),
    .B1(_05742_),
    .Y(_06114_));
 sky130_fd_sc_hd__a21o_1 _14579_ (.A1(_05928_),
    .A2(_06059_),
    .B1(_05742_),
    .X(_06125_));
 sky130_fd_sc_hd__o211a_1 _14580_ (.A1(net388),
    .A2(_06026_),
    .B1(_06092_),
    .C1(_06103_),
    .X(_06136_));
 sky130_fd_sc_hd__o2111a_1 _14581_ (.A1(net388),
    .A2(_06026_),
    .B1(net1),
    .C1(_06092_),
    .D1(_06103_),
    .X(_06147_));
 sky130_fd_sc_hd__o2111ai_4 _14582_ (.A1(net388),
    .A2(_06026_),
    .B1(net1),
    .C1(_06092_),
    .D1(_06103_),
    .Y(_06158_));
 sky130_fd_sc_hd__nor2_1 _14583_ (.A(net1),
    .B(_06136_),
    .Y(_06169_));
 sky130_fd_sc_hd__a211oi_1 _14584_ (.A1(_05687_),
    .A2(_05709_),
    .B1(_06147_),
    .C1(_06169_),
    .Y(_06180_));
 sky130_fd_sc_hd__a31o_1 _14585_ (.A1(_05687_),
    .A2(_05709_),
    .A3(_06136_),
    .B1(_06180_),
    .X(_06191_));
 sky130_fd_sc_hd__xnor2_1 _14586_ (.A(_05632_),
    .B(_06191_),
    .Y(net98));
 sky130_fd_sc_hd__and4bb_1 _14587_ (.A_N(_05272_),
    .B_N(_06191_),
    .C(_05611_),
    .D(_04613_),
    .X(_06212_));
 sky130_fd_sc_hd__nor4_4 _14588_ (.A(net12),
    .B(net1),
    .C(net23),
    .D(net26),
    .Y(_06223_));
 sky130_fd_sc_hd__nand3_4 _14589_ (.A(_05414_),
    .B(_03621_),
    .C(_03510_),
    .Y(_06234_));
 sky130_fd_sc_hd__a311oi_4 _14590_ (.A1(_03510_),
    .A2(_05414_),
    .A3(_03621_),
    .B1(_03399_),
    .C1(net27),
    .Y(_06245_));
 sky130_fd_sc_hd__nand3_4 _14591_ (.A(_06234_),
    .B(net25),
    .C(_03731_),
    .Y(_06256_));
 sky130_fd_sc_hd__a21oi_4 _14592_ (.A1(_06234_),
    .A2(net25),
    .B1(_03731_),
    .Y(_06267_));
 sky130_fd_sc_hd__o21ai_4 _14593_ (.A1(_03399_),
    .A2(_06223_),
    .B1(net27),
    .Y(_06278_));
 sky130_fd_sc_hd__a21oi_4 _14594_ (.A1(_06234_),
    .A2(net25),
    .B1(net27),
    .Y(_06289_));
 sky130_fd_sc_hd__o21bai_4 _14595_ (.A1(_03399_),
    .A2(_06223_),
    .B1_N(net27),
    .Y(_06300_));
 sky130_fd_sc_hd__o311a_4 _14596_ (.A1(net23),
    .A2(net26),
    .A3(_05425_),
    .B1(net27),
    .C1(net25),
    .X(_06310_));
 sky130_fd_sc_hd__nand3_4 _14597_ (.A(_06234_),
    .B(net27),
    .C(net25),
    .Y(_06321_));
 sky130_fd_sc_hd__nand2_8 _14598_ (.A(_06300_),
    .B(_06321_),
    .Y(_06332_));
 sky130_fd_sc_hd__nand2_8 _14599_ (.A(_06256_),
    .B(_06278_),
    .Y(_06343_));
 sky130_fd_sc_hd__a31oi_2 _14600_ (.A1(_06234_),
    .A2(net27),
    .A3(net25),
    .B1(_03178_),
    .Y(_06354_));
 sky130_fd_sc_hd__and3_1 _14601_ (.A(_06300_),
    .B(_06321_),
    .C(net33),
    .X(_06365_));
 sky130_fd_sc_hd__nand3_4 _14602_ (.A(_06300_),
    .B(_06321_),
    .C(net33),
    .Y(_06376_));
 sky130_fd_sc_hd__o2bb2ai_2 _14603_ (.A1_N(_05261_),
    .A2_N(_05950_),
    .B1(net386),
    .B2(_05873_),
    .Y(_06387_));
 sky130_fd_sc_hd__a21oi_1 _14604_ (.A1(_06256_),
    .A2(_06278_),
    .B1(_05873_),
    .Y(_06398_));
 sky130_fd_sc_hd__nand4_4 _14605_ (.A(_05862_),
    .B(_06300_),
    .C(_06321_),
    .D(net33),
    .Y(_06409_));
 sky130_fd_sc_hd__a21oi_1 _14606_ (.A1(_06354_),
    .A2(_06300_),
    .B1(_05862_),
    .Y(_06420_));
 sky130_fd_sc_hd__o2bb2ai_2 _14607_ (.A1_N(_06300_),
    .A2_N(_06354_),
    .B1(_05807_),
    .B2(_05829_),
    .Y(_06431_));
 sky130_fd_sc_hd__nand3_4 _14608_ (.A(_05895_),
    .B(_06387_),
    .C(_06431_),
    .Y(_06442_));
 sky130_fd_sc_hd__nand4_2 _14609_ (.A(_05895_),
    .B(_06387_),
    .C(_06409_),
    .D(_06431_),
    .Y(_06453_));
 sky130_fd_sc_hd__o2bb2ai_2 _14610_ (.A1_N(_05895_),
    .A2_N(_06387_),
    .B1(_06398_),
    .B2(_06420_),
    .Y(_06464_));
 sky130_fd_sc_hd__o221a_1 _14611_ (.A1(net408),
    .A2(_05152_),
    .B1(net393),
    .B2(net382),
    .C1(net33),
    .X(_06475_));
 sky130_fd_sc_hd__or4_2 _14612_ (.A(_03178_),
    .B(net404),
    .C(_06289_),
    .D(net391),
    .X(_06486_));
 sky130_fd_sc_hd__and3_1 _14613_ (.A(_06464_),
    .B(net404),
    .C(_06453_),
    .X(_06497_));
 sky130_fd_sc_hd__nand3_4 _14614_ (.A(_06464_),
    .B(net404),
    .C(_06453_),
    .Y(_06508_));
 sky130_fd_sc_hd__a31oi_1 _14615_ (.A1(_06464_),
    .A2(net404),
    .A3(_06453_),
    .B1(_06475_),
    .Y(_06519_));
 sky130_fd_sc_hd__a21oi_1 _14616_ (.A1(_06026_),
    .A2(net403),
    .B1(_06114_),
    .Y(_06530_));
 sky130_fd_sc_hd__o22ai_4 _14617_ (.A1(net398),
    .A2(net397),
    .B1(_06037_),
    .B2(_06114_),
    .Y(_06541_));
 sky130_fd_sc_hd__a31oi_4 _14618_ (.A1(_06048_),
    .A2(_06125_),
    .A3(net386),
    .B1(_05392_),
    .Y(_06552_));
 sky130_fd_sc_hd__o2111ai_4 _14619_ (.A1(net404),
    .A2(_06376_),
    .B1(_06508_),
    .C1(_06541_),
    .D1(_06552_),
    .Y(_06563_));
 sky130_fd_sc_hd__o2bb2ai_4 _14620_ (.A1_N(_06541_),
    .A2_N(_06552_),
    .B1(_06475_),
    .B2(_06497_),
    .Y(_06574_));
 sky130_fd_sc_hd__o21ai_1 _14621_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_06519_),
    .Y(_06585_));
 sky130_fd_sc_hd__a21oi_2 _14622_ (.A1(_06486_),
    .A2(_06508_),
    .B1(net386),
    .Y(_06596_));
 sky130_fd_sc_hd__and2_1 _14623_ (.A(_06563_),
    .B(_06574_),
    .X(_06607_));
 sky130_fd_sc_hd__or3_1 _14624_ (.A(net384),
    .B(net383),
    .C(_06607_),
    .X(_06617_));
 sky130_fd_sc_hd__a21oi_4 _14625_ (.A1(_06563_),
    .A2(_06574_),
    .B1(_05250_),
    .Y(_06628_));
 sky130_fd_sc_hd__a21o_1 _14626_ (.A1(_06563_),
    .A2(_06574_),
    .B1(_05250_),
    .X(_06639_));
 sky130_fd_sc_hd__and3_1 _14627_ (.A(_05250_),
    .B(_06563_),
    .C(_06574_),
    .X(_06650_));
 sky130_fd_sc_hd__nand3_1 _14628_ (.A(_05250_),
    .B(_06563_),
    .C(_06574_),
    .Y(_06661_));
 sky130_fd_sc_hd__a31oi_4 _14629_ (.A1(_05250_),
    .A2(_06563_),
    .A3(_06574_),
    .B1(_06158_),
    .Y(_06672_));
 sky130_fd_sc_hd__nand2_2 _14630_ (.A(_06661_),
    .B(_06147_),
    .Y(_06683_));
 sky130_fd_sc_hd__a21oi_1 _14631_ (.A1(_06639_),
    .A2(_06661_),
    .B1(_06147_),
    .Y(_06694_));
 sky130_fd_sc_hd__o21bai_1 _14632_ (.A1(_06628_),
    .A2(_06650_),
    .B1_N(_06147_),
    .Y(_06705_));
 sky130_fd_sc_hd__o21ai_1 _14633_ (.A1(_06628_),
    .A2(_06683_),
    .B1(net360),
    .Y(_06716_));
 sky130_fd_sc_hd__o221ai_4 _14634_ (.A1(net384),
    .A2(net383),
    .B1(_06628_),
    .B2(_06683_),
    .C1(_06705_),
    .Y(_06727_));
 sky130_fd_sc_hd__o22ai_1 _14635_ (.A1(net360),
    .A2(_06607_),
    .B1(_06694_),
    .B2(_06716_),
    .Y(_06738_));
 sky130_fd_sc_hd__a21oi_2 _14636_ (.A1(_06617_),
    .A2(_06727_),
    .B1(_03289_),
    .Y(_06749_));
 sky130_fd_sc_hd__nand2_1 _14637_ (.A(_06738_),
    .B(net1),
    .Y(_06760_));
 sky130_fd_sc_hd__o221a_1 _14638_ (.A1(net360),
    .A2(_06607_),
    .B1(_06694_),
    .B2(_06716_),
    .C1(_03289_),
    .X(_06771_));
 sky130_fd_sc_hd__o31ai_4 _14639_ (.A1(net55),
    .A2(net58),
    .A3(_05337_),
    .B1(net409),
    .Y(_06782_));
 sky130_fd_sc_hd__and2_4 _14640_ (.A(_06782_),
    .B(net59),
    .X(_06793_));
 sky130_fd_sc_hd__nand2_8 _14641_ (.A(_06782_),
    .B(net59),
    .Y(_06804_));
 sky130_fd_sc_hd__nor2_8 _14642_ (.A(net59),
    .B(_06782_),
    .Y(_06815_));
 sky130_fd_sc_hd__or2_4 _14643_ (.A(net59),
    .B(_06782_),
    .X(_06826_));
 sky130_fd_sc_hd__nand2_8 _14644_ (.A(_06804_),
    .B(_06826_),
    .Y(_06837_));
 sky130_fd_sc_hd__nor2_8 _14645_ (.A(net379),
    .B(net378),
    .Y(_06848_));
 sky130_fd_sc_hd__o22a_1 _14646_ (.A1(_06749_),
    .A2(_06771_),
    .B1(net379),
    .B2(net378),
    .X(_06859_));
 sky130_fd_sc_hd__a31o_1 _14647_ (.A1(_06617_),
    .A2(_06727_),
    .A3(_06848_),
    .B1(_06859_),
    .X(_06870_));
 sky130_fd_sc_hd__o21ai_1 _14648_ (.A1(_05051_),
    .A2(_06212_),
    .B1(_06870_),
    .Y(_06881_));
 sky130_fd_sc_hd__or3_1 _14649_ (.A(_05051_),
    .B(_06212_),
    .C(_06870_),
    .X(_06892_));
 sky130_fd_sc_hd__and2_1 _14650_ (.A(_06881_),
    .B(_06892_),
    .X(net109));
 sky130_fd_sc_hd__o2bb2a_1 _14651_ (.A1_N(_06212_),
    .A2_N(_06870_),
    .B1(_04832_),
    .B2(_04942_),
    .X(_06912_));
 sky130_fd_sc_hd__nand4_4 _14652_ (.A(_05414_),
    .B(_03731_),
    .C(_03621_),
    .D(_03510_),
    .Y(_06923_));
 sky130_fd_sc_hd__a31oi_1 _14653_ (.A1(_05753_),
    .A2(_03731_),
    .A3(_03621_),
    .B1(_03399_),
    .Y(_06934_));
 sky130_fd_sc_hd__and3_4 _14654_ (.A(_06923_),
    .B(net25),
    .C(_03841_),
    .X(_06945_));
 sky130_fd_sc_hd__a311o_4 _14655_ (.A1(_05753_),
    .A2(_03731_),
    .A3(_03621_),
    .B1(_03399_),
    .C1(net28),
    .X(_06956_));
 sky130_fd_sc_hd__a21oi_4 _14656_ (.A1(_06923_),
    .A2(net25),
    .B1(_03841_),
    .Y(_06967_));
 sky130_fd_sc_hd__a21o_4 _14657_ (.A1(_06923_),
    .A2(net25),
    .B1(_03841_),
    .X(_06978_));
 sky130_fd_sc_hd__and3_4 _14658_ (.A(_06923_),
    .B(net28),
    .C(net25),
    .X(_06989_));
 sky130_fd_sc_hd__o211ai_4 _14659_ (.A1(net27),
    .A2(_06234_),
    .B1(net28),
    .C1(net25),
    .Y(_07000_));
 sky130_fd_sc_hd__a21oi_4 _14660_ (.A1(_06923_),
    .A2(net25),
    .B1(net28),
    .Y(_07011_));
 sky130_fd_sc_hd__a21o_4 _14661_ (.A1(_06923_),
    .A2(net25),
    .B1(net28),
    .X(_07022_));
 sky130_fd_sc_hd__nand2_8 _14662_ (.A(net376),
    .B(_07022_),
    .Y(_07033_));
 sky130_fd_sc_hd__nand2_8 _14663_ (.A(_06956_),
    .B(_06978_),
    .Y(_07044_));
 sky130_fd_sc_hd__o21ai_1 _14664_ (.A1(net28),
    .A2(_06934_),
    .B1(net33),
    .Y(_07055_));
 sky130_fd_sc_hd__and3_1 _14665_ (.A(_07022_),
    .B(net33),
    .C(_07000_),
    .X(_07066_));
 sky130_fd_sc_hd__nand3_4 _14666_ (.A(_07022_),
    .B(net33),
    .C(_07000_),
    .Y(_07077_));
 sky130_fd_sc_hd__o221a_1 _14667_ (.A1(net408),
    .A2(_05152_),
    .B1(_06945_),
    .B2(net377),
    .C1(net33),
    .X(_07088_));
 sky130_fd_sc_hd__or4_1 _14668_ (.A(_03178_),
    .B(net404),
    .C(_06989_),
    .D(_07011_),
    .X(_07099_));
 sky130_fd_sc_hd__a21oi_2 _14669_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_06376_),
    .Y(_07110_));
 sky130_fd_sc_hd__a21o_1 _14670_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_06376_),
    .X(_07121_));
 sky130_fd_sc_hd__a31oi_2 _14671_ (.A1(_07000_),
    .A2(_07022_),
    .A3(net33),
    .B1(_06343_),
    .Y(_07132_));
 sky130_fd_sc_hd__o21ai_4 _14672_ (.A1(_06289_),
    .A2(net391),
    .B1(_07077_),
    .Y(_07143_));
 sky130_fd_sc_hd__o21ai_1 _14673_ (.A1(net393),
    .A2(net382),
    .B1(_07077_),
    .Y(_07154_));
 sky130_fd_sc_hd__o41ai_1 _14674_ (.A1(net393),
    .A2(net382),
    .A3(_06989_),
    .A4(_07055_),
    .B1(_07154_),
    .Y(_07165_));
 sky130_fd_sc_hd__o221ai_4 _14675_ (.A1(_05567_),
    .A2(_05851_),
    .B1(_05961_),
    .B2(_05884_),
    .C1(_06409_),
    .Y(_07176_));
 sky130_fd_sc_hd__o31a_2 _14676_ (.A1(_03178_),
    .A2(_05851_),
    .A3(_06332_),
    .B1(_06442_),
    .X(_07187_));
 sky130_fd_sc_hd__o2111ai_1 _14677_ (.A1(_06376_),
    .A2(_07033_),
    .B1(_07143_),
    .C1(_06409_),
    .D1(_06442_),
    .Y(_07198_));
 sky130_fd_sc_hd__o221ai_1 _14678_ (.A1(_05862_),
    .A2(_06365_),
    .B1(_07110_),
    .B2(_07132_),
    .C1(_07176_),
    .Y(_07209_));
 sky130_fd_sc_hd__o211ai_2 _14679_ (.A1(_05862_),
    .A2(_06365_),
    .B1(_07143_),
    .C1(_07176_),
    .Y(_07220_));
 sky130_fd_sc_hd__o211ai_2 _14680_ (.A1(_05862_),
    .A2(_06365_),
    .B1(_07176_),
    .C1(_07165_),
    .Y(_07231_));
 sky130_fd_sc_hd__o221ai_4 _14681_ (.A1(_05851_),
    .A2(_06376_),
    .B1(_07110_),
    .B2(_07132_),
    .C1(_06442_),
    .Y(_07241_));
 sky130_fd_sc_hd__a21oi_1 _14682_ (.A1(_07198_),
    .A2(_07209_),
    .B1(_05185_),
    .Y(_07252_));
 sky130_fd_sc_hd__nand3_2 _14683_ (.A(_07231_),
    .B(_07241_),
    .C(net404),
    .Y(_07263_));
 sky130_fd_sc_hd__o31a_1 _14684_ (.A1(_03178_),
    .A2(net404),
    .A3(_07033_),
    .B1(_07263_),
    .X(_07274_));
 sky130_fd_sc_hd__o21ai_1 _14685_ (.A1(net386),
    .A2(_06519_),
    .B1(_06530_),
    .Y(_07285_));
 sky130_fd_sc_hd__a32oi_4 _14686_ (.A1(_06508_),
    .A2(net386),
    .A3(_06486_),
    .B1(_06048_),
    .B2(_06125_),
    .Y(_07296_));
 sky130_fd_sc_hd__a311oi_1 _14687_ (.A1(_07231_),
    .A2(_07241_),
    .A3(net404),
    .B1(_05862_),
    .C1(_07088_),
    .Y(_07307_));
 sky130_fd_sc_hd__o221ai_4 _14688_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_07077_),
    .B2(net404),
    .C1(_07263_),
    .Y(_07318_));
 sky130_fd_sc_hd__a2bb2oi_1 _14689_ (.A1_N(_05763_),
    .A2_N(_05785_),
    .B1(_07099_),
    .B2(_07263_),
    .Y(_07329_));
 sky130_fd_sc_hd__o22ai_4 _14690_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_07088_),
    .B2(_07252_),
    .Y(_07340_));
 sky130_fd_sc_hd__o2bb2ai_1 _14691_ (.A1_N(_06585_),
    .A2_N(_07285_),
    .B1(_07307_),
    .B2(_07329_),
    .Y(_07351_));
 sky130_fd_sc_hd__o21ai_4 _14692_ (.A1(_06596_),
    .A2(_07296_),
    .B1(_07318_),
    .Y(_07362_));
 sky130_fd_sc_hd__o211ai_1 _14693_ (.A1(_06596_),
    .A2(_07296_),
    .B1(_07318_),
    .C1(_07340_),
    .Y(_07373_));
 sky130_fd_sc_hd__and3_1 _14694_ (.A(net388),
    .B(_07351_),
    .C(_07373_),
    .X(_07384_));
 sky130_fd_sc_hd__nand3_1 _14695_ (.A(net388),
    .B(_07351_),
    .C(_07373_),
    .Y(_07395_));
 sky130_fd_sc_hd__a211o_1 _14696_ (.A1(_07099_),
    .A2(_07263_),
    .B1(net402),
    .C1(net399),
    .X(_07406_));
 sky130_fd_sc_hd__inv_2 _14697_ (.A(_07406_),
    .Y(_07417_));
 sky130_fd_sc_hd__o31a_2 _14698_ (.A1(net402),
    .A2(net399),
    .A3(_07274_),
    .B1(_07395_),
    .X(_07428_));
 sky130_fd_sc_hd__nand3_4 _14699_ (.A(_06683_),
    .B(net386),
    .C(_06639_),
    .Y(_07439_));
 sky130_fd_sc_hd__o22ai_4 _14700_ (.A1(net398),
    .A2(net397),
    .B1(_06628_),
    .B2(_06672_),
    .Y(_07450_));
 sky130_fd_sc_hd__nand3_1 _14701_ (.A(_07450_),
    .B(net360),
    .C(_07439_),
    .Y(_07461_));
 sky130_fd_sc_hd__and4_1 _14702_ (.A(_07450_),
    .B(net360),
    .C(_07439_),
    .D(_07428_),
    .X(_07472_));
 sky130_fd_sc_hd__nand4_4 _14703_ (.A(_07450_),
    .B(net360),
    .C(_07439_),
    .D(_07428_),
    .Y(_07483_));
 sky130_fd_sc_hd__a31oi_2 _14704_ (.A1(_07450_),
    .A2(net360),
    .A3(_07439_),
    .B1(_07428_),
    .Y(_07494_));
 sky130_fd_sc_hd__o21ai_4 _14705_ (.A1(_07384_),
    .A2(_07417_),
    .B1(_07461_),
    .Y(_07505_));
 sky130_fd_sc_hd__nand3_1 _14706_ (.A(_07395_),
    .B(_07406_),
    .C(net386),
    .Y(_07516_));
 sky130_fd_sc_hd__a22o_1 _14707_ (.A1(_05458_),
    .A2(_05480_),
    .B1(_07395_),
    .B2(_07406_),
    .X(_07527_));
 sky130_fd_sc_hd__nor2_1 _14708_ (.A(_07472_),
    .B(_07494_),
    .Y(_07538_));
 sky130_fd_sc_hd__nand2_1 _14709_ (.A(_07483_),
    .B(_07505_),
    .Y(_07549_));
 sky130_fd_sc_hd__o211a_1 _14710_ (.A1(_05196_),
    .A2(_05218_),
    .B1(_07483_),
    .C1(_07505_),
    .X(_07559_));
 sky130_fd_sc_hd__o211ai_2 _14711_ (.A1(_05196_),
    .A2(_05218_),
    .B1(_07483_),
    .C1(_07505_),
    .Y(_07570_));
 sky130_fd_sc_hd__a21oi_2 _14712_ (.A1(_07483_),
    .A2(_07505_),
    .B1(_05250_),
    .Y(_07581_));
 sky130_fd_sc_hd__o21ai_2 _14713_ (.A1(_07472_),
    .A2(_07494_),
    .B1(net403),
    .Y(_07592_));
 sky130_fd_sc_hd__o21ai_2 _14714_ (.A1(_07559_),
    .A2(_07581_),
    .B1(_06760_),
    .Y(_07603_));
 sky130_fd_sc_hd__a31oi_2 _14715_ (.A1(_07592_),
    .A2(_06749_),
    .A3(_07570_),
    .B1(_06848_),
    .Y(_07614_));
 sky130_fd_sc_hd__a22oi_4 _14716_ (.A1(_06848_),
    .A2(_07549_),
    .B1(_07614_),
    .B2(_07603_),
    .Y(_07625_));
 sky130_fd_sc_hd__o2bb2ai_1 _14717_ (.A1_N(_07603_),
    .A2_N(_07614_),
    .B1(_06837_),
    .B2(_07538_),
    .Y(_07636_));
 sky130_fd_sc_hd__nor2_1 _14718_ (.A(_03289_),
    .B(_07625_),
    .Y(_07647_));
 sky130_fd_sc_hd__nand2_1 _14719_ (.A(_07636_),
    .B(net1),
    .Y(_07658_));
 sky130_fd_sc_hd__nor2_1 _14720_ (.A(net1),
    .B(_07636_),
    .Y(_07669_));
 sky130_fd_sc_hd__or4_4 _14721_ (.A(net55),
    .B(net58),
    .C(net59),
    .D(_05337_),
    .X(_07680_));
 sky130_fd_sc_hd__a21boi_4 _14722_ (.A1(_07680_),
    .A2(net409),
    .B1_N(net60),
    .Y(_07691_));
 sky130_fd_sc_hd__and3b_4 _14723_ (.A_N(net60),
    .B(_07680_),
    .C(net409),
    .X(_07702_));
 sky130_fd_sc_hd__or2_4 _14724_ (.A(net372),
    .B(net371),
    .X(_07713_));
 sky130_fd_sc_hd__nor2_8 _14725_ (.A(net372),
    .B(net371),
    .Y(_07724_));
 sky130_fd_sc_hd__or3_1 _14726_ (.A(_07625_),
    .B(net372),
    .C(net371),
    .X(_07735_));
 sky130_fd_sc_hd__o31a_1 _14727_ (.A1(_07724_),
    .A2(_07669_),
    .A3(_07647_),
    .B1(_07735_),
    .X(_07746_));
 sky130_fd_sc_hd__xnor2_1 _14728_ (.A(_06912_),
    .B(_07746_),
    .Y(net120));
 sky130_fd_sc_hd__and3_1 _14729_ (.A(_06212_),
    .B(_06870_),
    .C(_07746_),
    .X(_07767_));
 sky130_fd_sc_hd__nor2_4 _14730_ (.A(net27),
    .B(net28),
    .Y(_07778_));
 sky130_fd_sc_hd__nand4_4 _14731_ (.A(_05414_),
    .B(_07778_),
    .C(_03510_),
    .D(_03621_),
    .Y(_07789_));
 sky130_fd_sc_hd__a311oi_4 _14732_ (.A1(_05753_),
    .A2(_07778_),
    .A3(_03621_),
    .B1(net29),
    .C1(_03399_),
    .Y(_07800_));
 sky130_fd_sc_hd__a311o_4 _14733_ (.A1(_05753_),
    .A2(_07778_),
    .A3(_03621_),
    .B1(net29),
    .C1(_03399_),
    .X(_07811_));
 sky130_fd_sc_hd__a21oi_4 _14734_ (.A1(_07789_),
    .A2(net25),
    .B1(_03952_),
    .Y(_07822_));
 sky130_fd_sc_hd__a21o_4 _14735_ (.A1(_07789_),
    .A2(net25),
    .B1(_03952_),
    .X(_07833_));
 sky130_fd_sc_hd__a21oi_4 _14736_ (.A1(_07789_),
    .A2(net25),
    .B1(net29),
    .Y(_07844_));
 sky130_fd_sc_hd__a21o_4 _14737_ (.A1(_07789_),
    .A2(net410),
    .B1(net29),
    .X(_07855_));
 sky130_fd_sc_hd__o311a_4 _14738_ (.A1(net27),
    .A2(net28),
    .A3(_06234_),
    .B1(net29),
    .C1(net25),
    .X(_07866_));
 sky130_fd_sc_hd__a311o_4 _14739_ (.A1(_05753_),
    .A2(_07778_),
    .A3(_03621_),
    .B1(_03952_),
    .C1(_03399_),
    .X(_07877_));
 sky130_fd_sc_hd__nand2_8 _14740_ (.A(_07855_),
    .B(_07877_),
    .Y(_07888_));
 sky130_fd_sc_hd__nand2_8 _14741_ (.A(_07811_),
    .B(_07833_),
    .Y(_07899_));
 sky130_fd_sc_hd__a31o_1 _14742_ (.A1(_07789_),
    .A2(net29),
    .A3(net25),
    .B1(_03178_),
    .X(_07910_));
 sky130_fd_sc_hd__and3_1 _14743_ (.A(_07855_),
    .B(_07877_),
    .C(net33),
    .X(_07921_));
 sky130_fd_sc_hd__o21ai_4 _14744_ (.A1(net390),
    .A2(net370),
    .B1(net33),
    .Y(_07931_));
 sky130_fd_sc_hd__o22ai_4 _14745_ (.A1(net369),
    .A2(_07910_),
    .B1(_06989_),
    .B2(_07011_),
    .Y(_07942_));
 sky130_fd_sc_hd__and3_1 _14746_ (.A(_07044_),
    .B(_07899_),
    .C(net33),
    .X(_07953_));
 sky130_fd_sc_hd__o31a_2 _14747_ (.A1(net369),
    .A2(_07866_),
    .A3(_07077_),
    .B1(_07942_),
    .X(_07964_));
 sky130_fd_sc_hd__o21ai_1 _14748_ (.A1(_07077_),
    .A2(_07888_),
    .B1(_07942_),
    .Y(_07975_));
 sky130_fd_sc_hd__o211ai_4 _14749_ (.A1(_07077_),
    .A2(_06332_),
    .B1(_06409_),
    .C1(_06442_),
    .Y(_07986_));
 sky130_fd_sc_hd__o211ai_4 _14750_ (.A1(_06343_),
    .A2(_07066_),
    .B1(_07964_),
    .C1(_07986_),
    .Y(_07997_));
 sky130_fd_sc_hd__o211ai_4 _14751_ (.A1(_07077_),
    .A2(_06332_),
    .B1(_07975_),
    .C1(_07220_),
    .Y(_08008_));
 sky130_fd_sc_hd__nand3_1 _14752_ (.A(_07997_),
    .B(_08008_),
    .C(net404),
    .Y(_08019_));
 sky130_fd_sc_hd__o221a_2 _14753_ (.A1(net408),
    .A2(_05152_),
    .B1(net390),
    .B2(net370),
    .C1(net33),
    .X(_08030_));
 sky130_fd_sc_hd__or4_1 _14754_ (.A(_03178_),
    .B(net404),
    .C(net369),
    .D(_07866_),
    .X(_08041_));
 sky130_fd_sc_hd__a31oi_4 _14755_ (.A1(_07997_),
    .A2(_08008_),
    .A3(net404),
    .B1(_08030_),
    .Y(_08052_));
 sky130_fd_sc_hd__a31o_1 _14756_ (.A1(_07997_),
    .A2(_08008_),
    .A3(net404),
    .B1(_08030_),
    .X(_08063_));
 sky130_fd_sc_hd__a311o_2 _14757_ (.A1(_07997_),
    .A2(_08008_),
    .A3(net404),
    .B1(_08030_),
    .C1(net388),
    .X(_08074_));
 sky130_fd_sc_hd__a21oi_2 _14758_ (.A1(_08019_),
    .A2(_08041_),
    .B1(_06332_),
    .Y(_08085_));
 sky130_fd_sc_hd__a22o_2 _14759_ (.A1(_06256_),
    .A2(_06278_),
    .B1(_08019_),
    .B2(_08041_),
    .X(_08096_));
 sky130_fd_sc_hd__o311a_1 _14760_ (.A1(_03178_),
    .A2(net404),
    .A3(_07888_),
    .B1(_06332_),
    .C1(_08019_),
    .X(_08107_));
 sky130_fd_sc_hd__a311o_1 _14761_ (.A1(_07997_),
    .A2(_08008_),
    .A3(net404),
    .B1(_08030_),
    .C1(_06343_),
    .X(_08118_));
 sky130_fd_sc_hd__o2bb2ai_1 _14762_ (.A1_N(_07340_),
    .A2_N(_07362_),
    .B1(_08085_),
    .B2(_08107_),
    .Y(_08129_));
 sky130_fd_sc_hd__o2111ai_4 _14763_ (.A1(_05851_),
    .A2(_07274_),
    .B1(_07362_),
    .C1(_08096_),
    .D1(_08118_),
    .Y(_08140_));
 sky130_fd_sc_hd__o211ai_4 _14764_ (.A1(net402),
    .A2(net399),
    .B1(_08129_),
    .C1(_08140_),
    .Y(_08151_));
 sky130_fd_sc_hd__o221a_1 _14765_ (.A1(_05851_),
    .A2(_07274_),
    .B1(_08085_),
    .B2(_08107_),
    .C1(_07362_),
    .X(_08162_));
 sky130_fd_sc_hd__a22oi_2 _14766_ (.A1(_06332_),
    .A2(_08052_),
    .B1(_07362_),
    .B2(_07340_),
    .Y(_08173_));
 sky130_fd_sc_hd__o2bb2ai_4 _14767_ (.A1_N(_07340_),
    .A2_N(_07362_),
    .B1(_08063_),
    .B2(_06343_),
    .Y(_08184_));
 sky130_fd_sc_hd__o22ai_2 _14768_ (.A1(net402),
    .A2(net399),
    .B1(_08085_),
    .B2(_08184_),
    .Y(_08195_));
 sky130_fd_sc_hd__nand2_1 _14769_ (.A(_07450_),
    .B(_07428_),
    .Y(_08206_));
 sky130_fd_sc_hd__o21ai_2 _14770_ (.A1(_06628_),
    .A2(_06672_),
    .B1(_07516_),
    .Y(_08217_));
 sky130_fd_sc_hd__o21ai_1 _14771_ (.A1(net385),
    .A2(_07428_),
    .B1(_08217_),
    .Y(_08228_));
 sky130_fd_sc_hd__a21oi_4 _14772_ (.A1(_08074_),
    .A2(_08151_),
    .B1(_05862_),
    .Y(_08239_));
 sky130_fd_sc_hd__o221ai_4 _14773_ (.A1(net388),
    .A2(_08052_),
    .B1(_08162_),
    .B2(_08195_),
    .C1(_05851_),
    .Y(_08250_));
 sky130_fd_sc_hd__o211a_1 _14774_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_08074_),
    .C1(_08151_),
    .X(_08261_));
 sky130_fd_sc_hd__o211ai_4 _14775_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_08074_),
    .C1(_08151_),
    .Y(_08272_));
 sky130_fd_sc_hd__nand3_4 _14776_ (.A(_08228_),
    .B(_08250_),
    .C(_08272_),
    .Y(_08283_));
 sky130_fd_sc_hd__o2bb2ai_4 _14777_ (.A1_N(_07439_),
    .A2_N(_08206_),
    .B1(_08239_),
    .B2(_08261_),
    .Y(_08294_));
 sky130_fd_sc_hd__o211ai_4 _14778_ (.A1(net384),
    .A2(net383),
    .B1(_08283_),
    .C1(_08294_),
    .Y(_08304_));
 sky130_fd_sc_hd__and3_1 _14779_ (.A(_05731_),
    .B(_08074_),
    .C(_08151_),
    .X(_08315_));
 sky130_fd_sc_hd__inv_2 _14780_ (.A(_08315_),
    .Y(_08326_));
 sky130_fd_sc_hd__a31oi_4 _14781_ (.A1(_08294_),
    .A2(net360),
    .A3(_08283_),
    .B1(_08315_),
    .Y(_08337_));
 sky130_fd_sc_hd__a21oi_1 _14782_ (.A1(_07549_),
    .A2(net403),
    .B1(_06749_),
    .Y(_08348_));
 sky130_fd_sc_hd__a31oi_2 _14783_ (.A1(_05250_),
    .A2(_07483_),
    .A3(_07505_),
    .B1(_06760_),
    .Y(_08359_));
 sky130_fd_sc_hd__nand2_1 _14784_ (.A(_07570_),
    .B(_06749_),
    .Y(_08370_));
 sky130_fd_sc_hd__o21ai_2 _14785_ (.A1(_05250_),
    .A2(_07538_),
    .B1(_08370_),
    .Y(_08381_));
 sky130_fd_sc_hd__nand3_2 _14786_ (.A(_08370_),
    .B(net386),
    .C(_07592_),
    .Y(_08392_));
 sky130_fd_sc_hd__o22ai_2 _14787_ (.A1(net398),
    .A2(net397),
    .B1(_07581_),
    .B2(_08359_),
    .Y(_08403_));
 sky130_fd_sc_hd__and4_1 _14788_ (.A(_08403_),
    .B(_06837_),
    .C(_08392_),
    .D(_08337_),
    .X(_08414_));
 sky130_fd_sc_hd__nand4_2 _14789_ (.A(_08403_),
    .B(_06837_),
    .C(_08392_),
    .D(_08337_),
    .Y(_08425_));
 sky130_fd_sc_hd__a31oi_1 _14790_ (.A1(_08403_),
    .A2(_06837_),
    .A3(_08392_),
    .B1(_08337_),
    .Y(_08436_));
 sky130_fd_sc_hd__a31o_1 _14791_ (.A1(_08403_),
    .A2(_06837_),
    .A3(_08392_),
    .B1(_08337_),
    .X(_08447_));
 sky130_fd_sc_hd__a21oi_2 _14792_ (.A1(_08304_),
    .A2(_08326_),
    .B1(_06837_),
    .Y(_08458_));
 sky130_fd_sc_hd__a311oi_1 _14793_ (.A1(_08294_),
    .A2(net360),
    .A3(_08283_),
    .B1(_08315_),
    .C1(_05556_),
    .Y(_08469_));
 sky130_fd_sc_hd__nand3_2 _14794_ (.A(_08304_),
    .B(_08326_),
    .C(net385),
    .Y(_08480_));
 sky130_fd_sc_hd__a21oi_4 _14795_ (.A1(_08304_),
    .A2(_08326_),
    .B1(net385),
    .Y(_08491_));
 sky130_fd_sc_hd__a22o_1 _14796_ (.A1(_05458_),
    .A2(_05480_),
    .B1(_08304_),
    .B2(_08326_),
    .X(_08502_));
 sky130_fd_sc_hd__o211ai_2 _14797_ (.A1(net385),
    .A2(_08337_),
    .B1(_08480_),
    .C1(_08381_),
    .Y(_08513_));
 sky130_fd_sc_hd__o22ai_2 _14798_ (.A1(_07559_),
    .A2(_08348_),
    .B1(_08469_),
    .B2(_08491_),
    .Y(_08524_));
 sky130_fd_sc_hd__a31oi_4 _14799_ (.A1(_08524_),
    .A2(_06837_),
    .A3(_08513_),
    .B1(_08458_),
    .Y(_08535_));
 sky130_fd_sc_hd__a31o_1 _14800_ (.A1(_08524_),
    .A2(_06837_),
    .A3(_08513_),
    .B1(_08458_),
    .X(_08546_));
 sky130_fd_sc_hd__o211ai_2 _14801_ (.A1(_05196_),
    .A2(_05218_),
    .B1(_08425_),
    .C1(_08447_),
    .Y(_08557_));
 sky130_fd_sc_hd__a21oi_1 _14802_ (.A1(_08425_),
    .A2(_08447_),
    .B1(_05250_),
    .Y(_08568_));
 sky130_fd_sc_hd__o21ai_2 _14803_ (.A1(_08414_),
    .A2(_08436_),
    .B1(net403),
    .Y(_08579_));
 sky130_fd_sc_hd__o2bb2ai_1 _14804_ (.A1_N(_08557_),
    .A2_N(_08579_),
    .B1(_03289_),
    .B2(_07625_),
    .Y(_08590_));
 sky130_fd_sc_hd__a31oi_2 _14805_ (.A1(_08579_),
    .A2(_07647_),
    .A3(_08557_),
    .B1(_07724_),
    .Y(_08601_));
 sky130_fd_sc_hd__a22oi_1 _14806_ (.A1(_07724_),
    .A2(_08546_),
    .B1(_08601_),
    .B2(_08590_),
    .Y(_08612_));
 sky130_fd_sc_hd__o2bb2ai_2 _14807_ (.A1_N(_08590_),
    .A2_N(_08601_),
    .B1(_07713_),
    .B2(_08535_),
    .Y(_08623_));
 sky130_fd_sc_hd__nor2_1 _14808_ (.A(_03289_),
    .B(_08612_),
    .Y(_08634_));
 sky130_fd_sc_hd__nand2_1 _14809_ (.A(_08623_),
    .B(net1),
    .Y(_08645_));
 sky130_fd_sc_hd__nor2_1 _14810_ (.A(net1),
    .B(_08623_),
    .Y(_08656_));
 sky130_fd_sc_hd__o21ai_4 _14811_ (.A1(net60),
    .A2(_07680_),
    .B1(net409),
    .Y(_08667_));
 sky130_fd_sc_hd__nor2_8 _14812_ (.A(net61),
    .B(_08667_),
    .Y(_08678_));
 sky130_fd_sc_hd__or2_4 _14813_ (.A(net61),
    .B(_08667_),
    .X(_08689_));
 sky130_fd_sc_hd__and2_4 _14814_ (.A(_08667_),
    .B(net61),
    .X(_08700_));
 sky130_fd_sc_hd__nand2_8 _14815_ (.A(_08667_),
    .B(net61),
    .Y(_08711_));
 sky130_fd_sc_hd__nand2_8 _14816_ (.A(_08689_),
    .B(_08711_),
    .Y(_08721_));
 sky130_fd_sc_hd__nor2_8 _14817_ (.A(net353),
    .B(net352),
    .Y(_08732_));
 sky130_fd_sc_hd__or3_1 _14818_ (.A(_08612_),
    .B(net353),
    .C(net352),
    .X(_08743_));
 sky130_fd_sc_hd__o31a_2 _14819_ (.A1(_08634_),
    .A2(_08656_),
    .A3(_08732_),
    .B1(_08743_),
    .X(_08754_));
 sky130_fd_sc_hd__o21ai_1 _14820_ (.A1(_05051_),
    .A2(_07767_),
    .B1(_08754_),
    .Y(_08765_));
 sky130_fd_sc_hd__a311o_1 _14821_ (.A1(_06212_),
    .A2(_06870_),
    .A3(_07746_),
    .B1(_08754_),
    .C1(_05051_),
    .X(_08776_));
 sky130_fd_sc_hd__and2_1 _14822_ (.A(_08765_),
    .B(_08776_),
    .X(net125));
 sky130_fd_sc_hd__o2bb2a_1 _14823_ (.A1_N(_07767_),
    .A2_N(_08754_),
    .B1(_04832_),
    .B2(_04942_),
    .X(_08797_));
 sky130_fd_sc_hd__nand4_4 _14824_ (.A(_05753_),
    .B(_07778_),
    .C(_03621_),
    .D(_03952_),
    .Y(_08808_));
 sky130_fd_sc_hd__o311a_4 _14825_ (.A1(net28),
    .A2(net29),
    .A3(_06923_),
    .B1(_04062_),
    .C1(net25),
    .X(_08819_));
 sky130_fd_sc_hd__a311o_4 _14826_ (.A1(_06223_),
    .A2(_07778_),
    .A3(_03952_),
    .B1(net30),
    .C1(_03399_),
    .X(_08830_));
 sky130_fd_sc_hd__a21oi_4 _14827_ (.A1(_08808_),
    .A2(net25),
    .B1(_04062_),
    .Y(_08841_));
 sky130_fd_sc_hd__a21o_4 _14828_ (.A1(_08808_),
    .A2(net410),
    .B1(_04062_),
    .X(_08852_));
 sky130_fd_sc_hd__o311a_4 _14829_ (.A1(net28),
    .A2(net29),
    .A3(_06923_),
    .B1(net30),
    .C1(net25),
    .X(_08863_));
 sky130_fd_sc_hd__o211ai_4 _14830_ (.A1(net29),
    .A2(_07789_),
    .B1(net30),
    .C1(net410),
    .Y(_08874_));
 sky130_fd_sc_hd__a21oi_4 _14831_ (.A1(_08808_),
    .A2(net410),
    .B1(net30),
    .Y(_08885_));
 sky130_fd_sc_hd__a21o_4 _14832_ (.A1(_08808_),
    .A2(net410),
    .B1(net30),
    .X(_08896_));
 sky130_fd_sc_hd__nand2_8 _14833_ (.A(_08874_),
    .B(_08896_),
    .Y(_08907_));
 sky130_fd_sc_hd__nand2_8 _14834_ (.A(_08830_),
    .B(_08852_),
    .Y(_08918_));
 sky130_fd_sc_hd__nand3_4 _14835_ (.A(_08896_),
    .B(net33),
    .C(_08874_),
    .Y(_08929_));
 sky130_fd_sc_hd__o21ai_1 _14836_ (.A1(net369),
    .A2(_07866_),
    .B1(_08929_),
    .Y(_08940_));
 sky130_fd_sc_hd__o21ai_4 _14837_ (.A1(_07931_),
    .A2(_08907_),
    .B1(_08940_),
    .Y(_08951_));
 sky130_fd_sc_hd__inv_2 _14838_ (.A(_08951_),
    .Y(_08962_));
 sky130_fd_sc_hd__a31oi_4 _14839_ (.A1(_07143_),
    .A2(_07986_),
    .A3(_07964_),
    .B1(_07953_),
    .Y(_08973_));
 sky130_fd_sc_hd__o21ai_1 _14840_ (.A1(_07033_),
    .A2(_07931_),
    .B1(_07997_),
    .Y(_08984_));
 sky130_fd_sc_hd__o211ai_4 _14841_ (.A1(_07888_),
    .A2(_07077_),
    .B1(_08951_),
    .C1(_07997_),
    .Y(_08995_));
 sky130_fd_sc_hd__nand2_2 _14842_ (.A(_08984_),
    .B(_08962_),
    .Y(_09006_));
 sky130_fd_sc_hd__o2111ai_4 _14843_ (.A1(_08951_),
    .A2(_08973_),
    .B1(_08995_),
    .C1(_05163_),
    .D1(_05141_),
    .Y(_09017_));
 sky130_fd_sc_hd__o221a_2 _14844_ (.A1(net408),
    .A2(_05152_),
    .B1(_08819_),
    .B2(net367),
    .C1(net33),
    .X(_09028_));
 sky130_fd_sc_hd__or4_1 _14845_ (.A(_03178_),
    .B(net404),
    .C(_08863_),
    .D(net366),
    .X(_09039_));
 sky130_fd_sc_hd__a31oi_4 _14846_ (.A1(_09006_),
    .A2(net404),
    .A3(_08995_),
    .B1(_09028_),
    .Y(_09050_));
 sky130_fd_sc_hd__a31o_2 _14847_ (.A1(_09006_),
    .A2(net404),
    .A3(_08995_),
    .B1(_09028_),
    .X(_09061_));
 sky130_fd_sc_hd__o311a_1 _14848_ (.A1(_03178_),
    .A2(net404),
    .A3(_08907_),
    .B1(_05392_),
    .C1(_09017_),
    .X(_09072_));
 sky130_fd_sc_hd__a311oi_2 _14849_ (.A1(_09006_),
    .A2(net404),
    .A3(_08995_),
    .B1(_09028_),
    .C1(_07044_),
    .Y(_09083_));
 sky130_fd_sc_hd__a311o_2 _14850_ (.A1(_09006_),
    .A2(net404),
    .A3(_08995_),
    .B1(_09028_),
    .C1(_07044_),
    .X(_09094_));
 sky130_fd_sc_hd__a21oi_1 _14851_ (.A1(_09017_),
    .A2(_09039_),
    .B1(_07033_),
    .Y(_09105_));
 sky130_fd_sc_hd__a22o_1 _14852_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_09017_),
    .B2(_09039_),
    .X(_09116_));
 sky130_fd_sc_hd__o221ai_2 _14853_ (.A1(_06332_),
    .A2(_08052_),
    .B1(_09083_),
    .B2(_09105_),
    .C1(_08184_),
    .Y(_09127_));
 sky130_fd_sc_hd__o211ai_1 _14854_ (.A1(_08085_),
    .A2(_08173_),
    .B1(_09094_),
    .C1(_09116_),
    .Y(_09137_));
 sky130_fd_sc_hd__o2111ai_4 _14855_ (.A1(_06332_),
    .A2(_08052_),
    .B1(_08184_),
    .C1(_09094_),
    .D1(_09116_),
    .Y(_09148_));
 sky130_fd_sc_hd__o22ai_2 _14856_ (.A1(_08085_),
    .A2(_08173_),
    .B1(_09083_),
    .B2(_09105_),
    .Y(_09159_));
 sky130_fd_sc_hd__o211ai_2 _14857_ (.A1(net402),
    .A2(net399),
    .B1(_09148_),
    .C1(_09159_),
    .Y(_09170_));
 sky130_fd_sc_hd__or3_1 _14858_ (.A(net402),
    .B(net399),
    .C(_09050_),
    .X(_09181_));
 sky130_fd_sc_hd__nand3_1 _14859_ (.A(net388),
    .B(_09127_),
    .C(_09137_),
    .Y(_09192_));
 sky130_fd_sc_hd__a311oi_1 _14860_ (.A1(net388),
    .A2(_09148_),
    .A3(_09159_),
    .B1(_06332_),
    .C1(_09072_),
    .Y(_09203_));
 sky130_fd_sc_hd__o211ai_4 _14861_ (.A1(net388),
    .A2(_09061_),
    .B1(_09170_),
    .C1(_06343_),
    .Y(_09214_));
 sky130_fd_sc_hd__a31oi_1 _14862_ (.A1(net388),
    .A2(_09127_),
    .A3(_09137_),
    .B1(_06343_),
    .Y(_09225_));
 sky130_fd_sc_hd__o221ai_4 _14863_ (.A1(_06289_),
    .A2(net391),
    .B1(_09050_),
    .B2(net388),
    .C1(_09192_),
    .Y(_09236_));
 sky130_fd_sc_hd__o211a_1 _14864_ (.A1(net385),
    .A2(_07428_),
    .B1(_08217_),
    .C1(_08272_),
    .X(_09247_));
 sky130_fd_sc_hd__o211ai_1 _14865_ (.A1(net385),
    .A2(_07428_),
    .B1(_08217_),
    .C1(_08272_),
    .Y(_09258_));
 sky130_fd_sc_hd__a31oi_4 _14866_ (.A1(_07527_),
    .A2(_08217_),
    .A3(_08272_),
    .B1(_08239_),
    .Y(_09269_));
 sky130_fd_sc_hd__nand2_1 _14867_ (.A(_08250_),
    .B(_09258_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand3_4 _14868_ (.A(_09269_),
    .B(_09236_),
    .C(_09214_),
    .Y(_09291_));
 sky130_fd_sc_hd__o2bb2ai_4 _14869_ (.A1_N(_09214_),
    .A2_N(_09236_),
    .B1(_09247_),
    .B2(_08239_),
    .Y(_09302_));
 sky130_fd_sc_hd__o211ai_2 _14870_ (.A1(net384),
    .A2(net383),
    .B1(_09291_),
    .C1(_09302_),
    .Y(_09313_));
 sky130_fd_sc_hd__o311a_2 _14871_ (.A1(net402),
    .A2(_09061_),
    .A3(net399),
    .B1(_05731_),
    .C1(_09170_),
    .X(_09324_));
 sky130_fd_sc_hd__a311o_1 _14872_ (.A1(net388),
    .A2(_09148_),
    .A3(_09159_),
    .B1(net360),
    .C1(_09072_),
    .X(_09335_));
 sky130_fd_sc_hd__a31oi_4 _14873_ (.A1(_09302_),
    .A2(net360),
    .A3(_09291_),
    .B1(_09324_),
    .Y(_09346_));
 sky130_fd_sc_hd__o21ai_1 _14874_ (.A1(_07581_),
    .A2(_08359_),
    .B1(_08480_),
    .Y(_09357_));
 sky130_fd_sc_hd__a22oi_2 _14875_ (.A1(_07592_),
    .A2(_08370_),
    .B1(_08337_),
    .B2(net386),
    .Y(_09368_));
 sky130_fd_sc_hd__a21oi_4 _14876_ (.A1(_08381_),
    .A2(_08480_),
    .B1(_08491_),
    .Y(_09379_));
 sky130_fd_sc_hd__a311oi_4 _14877_ (.A1(_09302_),
    .A2(net360),
    .A3(_09291_),
    .B1(_09324_),
    .C1(_05862_),
    .Y(_09390_));
 sky130_fd_sc_hd__a311o_1 _14878_ (.A1(_09302_),
    .A2(net360),
    .A3(_09291_),
    .B1(_09324_),
    .C1(_05862_),
    .X(_09401_));
 sky130_fd_sc_hd__a21oi_1 _14879_ (.A1(_09313_),
    .A2(_09335_),
    .B1(_05851_),
    .Y(_09412_));
 sky130_fd_sc_hd__a22o_1 _14880_ (.A1(_05774_),
    .A2(_05796_),
    .B1(_09313_),
    .B2(_09335_),
    .X(_09423_));
 sky130_fd_sc_hd__o221ai_4 _14881_ (.A1(_05851_),
    .A2(_09346_),
    .B1(_08491_),
    .B2(_09368_),
    .C1(_09401_),
    .Y(_09434_));
 sky130_fd_sc_hd__o21ai_2 _14882_ (.A1(_09390_),
    .A2(_09412_),
    .B1(_09379_),
    .Y(_09445_));
 sky130_fd_sc_hd__o211ai_2 _14883_ (.A1(net379),
    .A2(net378),
    .B1(_09434_),
    .C1(_09445_),
    .Y(_09456_));
 sky130_fd_sc_hd__a21oi_1 _14884_ (.A1(_09313_),
    .A2(_09335_),
    .B1(_06837_),
    .Y(_09467_));
 sky130_fd_sc_hd__or3_1 _14885_ (.A(net379),
    .B(net378),
    .C(_09346_),
    .X(_09478_));
 sky130_fd_sc_hd__a31oi_4 _14886_ (.A1(_09434_),
    .A2(_09445_),
    .A3(_06837_),
    .B1(_09467_),
    .Y(_09489_));
 sky130_fd_sc_hd__o22ai_2 _14887_ (.A1(_03289_),
    .A2(_07625_),
    .B1(_05250_),
    .B2(_08535_),
    .Y(_09500_));
 sky130_fd_sc_hd__a31oi_1 _14888_ (.A1(_05250_),
    .A2(_08425_),
    .A3(_08447_),
    .B1(_07658_),
    .Y(_09511_));
 sky130_fd_sc_hd__nand2_2 _14889_ (.A(_08557_),
    .B(_07647_),
    .Y(_09522_));
 sky130_fd_sc_hd__o21ai_1 _14890_ (.A1(_05250_),
    .A2(_08535_),
    .B1(_09522_),
    .Y(_09533_));
 sky130_fd_sc_hd__o31a_1 _14891_ (.A1(_05196_),
    .A2(_05218_),
    .A3(_08535_),
    .B1(_09522_),
    .X(_09544_));
 sky130_fd_sc_hd__o211ai_4 _14892_ (.A1(_08546_),
    .A2(net403),
    .B1(_05556_),
    .C1(_09500_),
    .Y(_09555_));
 sky130_fd_sc_hd__o221ai_4 _14893_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_08535_),
    .B2(_05250_),
    .C1(_09522_),
    .Y(_09566_));
 sky130_fd_sc_hd__and4_1 _14894_ (.A(_09555_),
    .B(_09566_),
    .C(_07713_),
    .D(_09489_),
    .X(_09576_));
 sky130_fd_sc_hd__nand4_4 _14895_ (.A(_09555_),
    .B(_09566_),
    .C(_07713_),
    .D(_09489_),
    .Y(_09587_));
 sky130_fd_sc_hd__a31oi_2 _14896_ (.A1(_09555_),
    .A2(_09566_),
    .A3(_07713_),
    .B1(_09489_),
    .Y(_09598_));
 sky130_fd_sc_hd__a31o_2 _14897_ (.A1(_09555_),
    .A2(_09566_),
    .A3(_07713_),
    .B1(_09489_),
    .X(_09609_));
 sky130_fd_sc_hd__o311a_1 _14898_ (.A1(net379),
    .A2(net378),
    .A3(_09346_),
    .B1(net385),
    .C1(_09456_),
    .X(_09620_));
 sky130_fd_sc_hd__nand3_1 _14899_ (.A(_09456_),
    .B(_09478_),
    .C(net385),
    .Y(_09631_));
 sky130_fd_sc_hd__a21oi_1 _14900_ (.A1(_09456_),
    .A2(_09478_),
    .B1(net385),
    .Y(_09642_));
 sky130_fd_sc_hd__a22o_1 _14901_ (.A1(_05458_),
    .A2(_05480_),
    .B1(_09456_),
    .B2(_09478_),
    .X(_09653_));
 sky130_fd_sc_hd__o211a_1 _14902_ (.A1(_09576_),
    .A2(_09598_),
    .B1(_08689_),
    .C1(_08711_),
    .X(_09664_));
 sky130_fd_sc_hd__o211ai_2 _14903_ (.A1(_05196_),
    .A2(_05218_),
    .B1(_09587_),
    .C1(_09609_),
    .Y(_09675_));
 sky130_fd_sc_hd__a21oi_2 _14904_ (.A1(_09587_),
    .A2(_09609_),
    .B1(_05250_),
    .Y(_09686_));
 sky130_fd_sc_hd__o21ai_2 _14905_ (.A1(_09576_),
    .A2(_09598_),
    .B1(net403),
    .Y(_09697_));
 sky130_fd_sc_hd__a22o_1 _14906_ (.A1(_08623_),
    .A2(net1),
    .B1(_09697_),
    .B2(_09675_),
    .X(_09708_));
 sky130_fd_sc_hd__nand4_1 _14907_ (.A(_08623_),
    .B(_09675_),
    .C(_09697_),
    .D(net1),
    .Y(_09719_));
 sky130_fd_sc_hd__a31oi_2 _14908_ (.A1(_09708_),
    .A2(_09719_),
    .A3(_08721_),
    .B1(_09664_),
    .Y(_09730_));
 sky130_fd_sc_hd__a31o_1 _14909_ (.A1(_09708_),
    .A2(_09719_),
    .A3(_08721_),
    .B1(_09664_),
    .X(_09741_));
 sky130_fd_sc_hd__or3_4 _14910_ (.A(net60),
    .B(net61),
    .C(_07680_),
    .X(_09752_));
 sky130_fd_sc_hd__o311a_4 _14911_ (.A1(net60),
    .A2(net61),
    .A3(_07680_),
    .B1(net62),
    .C1(net409),
    .X(_09763_));
 sky130_fd_sc_hd__a21oi_4 _14912_ (.A1(_09752_),
    .A2(net409),
    .B1(net62),
    .Y(_09774_));
 sky130_fd_sc_hd__a21boi_4 _14913_ (.A1(_09752_),
    .A2(net409),
    .B1_N(net62),
    .Y(_09785_));
 sky130_fd_sc_hd__clkinv_4 _14914_ (.A(net350),
    .Y(_09796_));
 sky130_fd_sc_hd__and3b_4 _14915_ (.A_N(net62),
    .B(_09752_),
    .C(net409),
    .X(_09807_));
 sky130_fd_sc_hd__clkinv_4 _14916_ (.A(net349),
    .Y(_09818_));
 sky130_fd_sc_hd__nor2_8 _14917_ (.A(_09763_),
    .B(_09774_),
    .Y(_09829_));
 sky130_fd_sc_hd__nor2_8 _14918_ (.A(net350),
    .B(net349),
    .Y(_09840_));
 sky130_fd_sc_hd__o21ai_1 _14919_ (.A1(_03289_),
    .A2(_09840_),
    .B1(_09741_),
    .Y(_09851_));
 sky130_fd_sc_hd__nand2_1 _14920_ (.A(_09741_),
    .B(net1),
    .Y(_09862_));
 sky130_fd_sc_hd__o31a_1 _14921_ (.A1(_03289_),
    .A2(_09741_),
    .A3(_09840_),
    .B1(_09851_),
    .X(_09873_));
 sky130_fd_sc_hd__xnor2_1 _14922_ (.A(_08797_),
    .B(_09873_),
    .Y(net126));
 sky130_fd_sc_hd__nand3_2 _14923_ (.A(_07767_),
    .B(_08754_),
    .C(_09873_),
    .Y(_09894_));
 sky130_fd_sc_hd__and4_2 _14924_ (.A(_06223_),
    .B(_07778_),
    .C(_03952_),
    .D(_04062_),
    .X(_09905_));
 sky130_fd_sc_hd__nand4_4 _14925_ (.A(_06223_),
    .B(_07778_),
    .C(_03952_),
    .D(_04062_),
    .Y(_09916_));
 sky130_fd_sc_hd__and3b_4 _14926_ (.A_N(net31),
    .B(_09916_),
    .C(net410),
    .X(_09927_));
 sky130_fd_sc_hd__or3_4 _14927_ (.A(_03399_),
    .B(net31),
    .C(_09905_),
    .X(_09938_));
 sky130_fd_sc_hd__o21a_4 _14928_ (.A1(_03399_),
    .A2(_09905_),
    .B1(net31),
    .X(_09949_));
 sky130_fd_sc_hd__o21ai_4 _14929_ (.A1(_03399_),
    .A2(_09905_),
    .B1(net31),
    .Y(_09960_));
 sky130_fd_sc_hd__o311a_4 _14930_ (.A1(net29),
    .A2(net30),
    .A3(_07789_),
    .B1(net31),
    .C1(net25),
    .X(_09971_));
 sky130_fd_sc_hd__o211ai_4 _14931_ (.A1(net30),
    .A2(_08808_),
    .B1(net31),
    .C1(net410),
    .Y(_09982_));
 sky130_fd_sc_hd__a21oi_4 _14932_ (.A1(_09916_),
    .A2(net25),
    .B1(net31),
    .Y(_09993_));
 sky130_fd_sc_hd__a21o_4 _14933_ (.A1(_09916_),
    .A2(net410),
    .B1(net31),
    .X(_10004_));
 sky130_fd_sc_hd__nand2_8 _14934_ (.A(_09982_),
    .B(_10004_),
    .Y(_10015_));
 sky130_fd_sc_hd__nor2_8 _14935_ (.A(net365),
    .B(net362),
    .Y(_10025_));
 sky130_fd_sc_hd__or3_4 _14936_ (.A(_03178_),
    .B(_09971_),
    .C(_09993_),
    .X(_10036_));
 sky130_fd_sc_hd__o32a_1 _14937_ (.A1(_03178_),
    .A2(_09971_),
    .A3(net363),
    .B1(net408),
    .B2(_05152_),
    .X(_10047_));
 sky130_fd_sc_hd__a22oi_1 _14938_ (.A1(_07921_),
    .A2(_08918_),
    .B1(_08984_),
    .B2(_08962_),
    .Y(_10058_));
 sky130_fd_sc_hd__o22ai_4 _14939_ (.A1(_07931_),
    .A2(_08907_),
    .B1(_08951_),
    .B2(_08973_),
    .Y(_10069_));
 sky130_fd_sc_hd__a31o_2 _14940_ (.A1(net33),
    .A2(_09982_),
    .A3(_10004_),
    .B1(_08918_),
    .X(_10080_));
 sky130_fd_sc_hd__and3_1 _14941_ (.A(net348),
    .B(_08907_),
    .C(net33),
    .X(_10091_));
 sky130_fd_sc_hd__o32a_1 _14942_ (.A1(_03178_),
    .A2(_09971_),
    .A3(net363),
    .B1(_08819_),
    .B2(net367),
    .X(_10102_));
 sky130_fd_sc_hd__o31a_1 _14943_ (.A1(_08929_),
    .A2(_09971_),
    .A3(net363),
    .B1(_10080_),
    .X(_10113_));
 sky130_fd_sc_hd__o21ai_2 _14944_ (.A1(_08929_),
    .A2(_10015_),
    .B1(_10080_),
    .Y(_10124_));
 sky130_fd_sc_hd__o221ai_4 _14945_ (.A1(_07931_),
    .A2(_08907_),
    .B1(_08951_),
    .B2(_08973_),
    .C1(_10124_),
    .Y(_10135_));
 sky130_fd_sc_hd__o21ai_4 _14946_ (.A1(_10091_),
    .A2(_10102_),
    .B1(_10069_),
    .Y(_10146_));
 sky130_fd_sc_hd__a21oi_1 _14947_ (.A1(_10135_),
    .A2(_10146_),
    .B1(_05185_),
    .Y(_10157_));
 sky130_fd_sc_hd__and3_1 _14948_ (.A(net348),
    .B(net33),
    .C(_05185_),
    .X(_10168_));
 sky130_fd_sc_hd__or4_1 _14949_ (.A(_03178_),
    .B(net404),
    .C(_09971_),
    .D(net363),
    .X(_10179_));
 sky130_fd_sc_hd__nand3_2 _14950_ (.A(_10146_),
    .B(net404),
    .C(_10135_),
    .Y(_10190_));
 sky130_fd_sc_hd__a31oi_4 _14951_ (.A1(_10146_),
    .A2(net404),
    .A3(_10135_),
    .B1(_10168_),
    .Y(_10201_));
 sky130_fd_sc_hd__a21oi_2 _14952_ (.A1(_10179_),
    .A2(_10190_),
    .B1(net388),
    .Y(_10212_));
 sky130_fd_sc_hd__inv_2 _14953_ (.A(_10212_),
    .Y(_10223_));
 sky130_fd_sc_hd__o311a_1 _14954_ (.A1(_03178_),
    .A2(net404),
    .A3(_10015_),
    .B1(_07888_),
    .C1(_10190_),
    .X(_10234_));
 sky130_fd_sc_hd__o21ai_2 _14955_ (.A1(net369),
    .A2(_07866_),
    .B1(_10201_),
    .Y(_10245_));
 sky130_fd_sc_hd__a21oi_2 _14956_ (.A1(_10179_),
    .A2(_10190_),
    .B1(_07888_),
    .Y(_10256_));
 sky130_fd_sc_hd__o211ai_4 _14957_ (.A1(_07033_),
    .A2(_09050_),
    .B1(_08184_),
    .C1(_08096_),
    .Y(_10267_));
 sky130_fd_sc_hd__o21ai_1 _14958_ (.A1(_07044_),
    .A2(_09061_),
    .B1(_10267_),
    .Y(_10278_));
 sky130_fd_sc_hd__o21ai_1 _14959_ (.A1(_10234_),
    .A2(_10256_),
    .B1(_10278_),
    .Y(_10289_));
 sky130_fd_sc_hd__o221ai_4 _14960_ (.A1(_07044_),
    .A2(_09061_),
    .B1(_07888_),
    .B2(_10201_),
    .C1(_10267_),
    .Y(_10300_));
 sky130_fd_sc_hd__o211ai_4 _14961_ (.A1(_10300_),
    .A2(_10234_),
    .B1(net388),
    .C1(_10289_),
    .Y(_10311_));
 sky130_fd_sc_hd__o31a_1 _14962_ (.A1(net388),
    .A2(_10047_),
    .A3(_10157_),
    .B1(_10311_),
    .X(_10322_));
 sky130_fd_sc_hd__or4b_2 _14963_ (.A(net384),
    .B(net383),
    .C(_10212_),
    .D_N(_10311_),
    .X(_10333_));
 sky130_fd_sc_hd__o21ai_1 _14964_ (.A1(_06989_),
    .A2(_07011_),
    .B1(_10311_),
    .Y(_10344_));
 sky130_fd_sc_hd__o311a_4 _14965_ (.A1(net388),
    .A2(_10047_),
    .A3(_10157_),
    .B1(_07033_),
    .C1(_10311_),
    .X(_10355_));
 sky130_fd_sc_hd__a2bb2oi_1 _14966_ (.A1_N(_06945_),
    .A2_N(net377),
    .B1(_10223_),
    .B2(_10311_),
    .Y(_10366_));
 sky130_fd_sc_hd__a22o_1 _14967_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_10223_),
    .B2(_10311_),
    .X(_10377_));
 sky130_fd_sc_hd__a22oi_2 _14968_ (.A1(_09181_),
    .A2(_09225_),
    .B1(_09280_),
    .B2(_09214_),
    .Y(_10388_));
 sky130_fd_sc_hd__o21ai_2 _14969_ (.A1(_09203_),
    .A2(_09269_),
    .B1(_09236_),
    .Y(_10399_));
 sky130_fd_sc_hd__o211ai_1 _14970_ (.A1(_10344_),
    .A2(_10212_),
    .B1(_10399_),
    .C1(_10377_),
    .Y(_10410_));
 sky130_fd_sc_hd__o21ai_1 _14971_ (.A1(_10355_),
    .A2(_10366_),
    .B1(_10388_),
    .Y(_10421_));
 sky130_fd_sc_hd__nand3_2 _14972_ (.A(_10421_),
    .B(net360),
    .C(_10410_),
    .Y(_10432_));
 sky130_fd_sc_hd__or3_1 _14973_ (.A(net384),
    .B(net383),
    .C(_10322_),
    .X(_10443_));
 sky130_fd_sc_hd__o21ai_1 _14974_ (.A1(_10355_),
    .A2(_10366_),
    .B1(_10399_),
    .Y(_10454_));
 sky130_fd_sc_hd__o211ai_1 _14975_ (.A1(_10212_),
    .A2(_10344_),
    .B1(_10388_),
    .C1(_10377_),
    .Y(_10465_));
 sky130_fd_sc_hd__nand3_2 _14976_ (.A(_10454_),
    .B(_10465_),
    .C(net360),
    .Y(_10476_));
 sky130_fd_sc_hd__and3_4 _14977_ (.A(_06848_),
    .B(_10333_),
    .C(_10432_),
    .X(_10486_));
 sky130_fd_sc_hd__a211o_1 _14978_ (.A1(_10443_),
    .A2(_10476_),
    .B1(net379),
    .C1(net378),
    .X(_10497_));
 sky130_fd_sc_hd__a2bb2oi_2 _14979_ (.A1_N(net393),
    .A2_N(net382),
    .B1(_10443_),
    .B2(_10476_),
    .Y(_10508_));
 sky130_fd_sc_hd__o211ai_4 _14980_ (.A1(net393),
    .A2(net382),
    .B1(_10333_),
    .C1(_10432_),
    .Y(_10519_));
 sky130_fd_sc_hd__o221ai_4 _14981_ (.A1(net380),
    .A2(net391),
    .B1(_10322_),
    .B2(net360),
    .C1(_10476_),
    .Y(_10530_));
 sky130_fd_sc_hd__inv_2 _14982_ (.A(_10530_),
    .Y(_10541_));
 sky130_fd_sc_hd__o211a_1 _14983_ (.A1(_05851_),
    .A2(_09346_),
    .B1(_09357_),
    .C1(_08502_),
    .X(_10552_));
 sky130_fd_sc_hd__a21oi_1 _14984_ (.A1(_08502_),
    .A2(_09357_),
    .B1(_09390_),
    .Y(_10563_));
 sky130_fd_sc_hd__o21ai_4 _14985_ (.A1(_09390_),
    .A2(_09379_),
    .B1(_09423_),
    .Y(_10574_));
 sky130_fd_sc_hd__o2bb2ai_1 _14986_ (.A1_N(_10519_),
    .A2_N(_10530_),
    .B1(_10563_),
    .B2(_09412_),
    .Y(_10585_));
 sky130_fd_sc_hd__o2111ai_1 _14987_ (.A1(_09379_),
    .A2(_09390_),
    .B1(_09423_),
    .C1(_10519_),
    .D1(_10530_),
    .Y(_10596_));
 sky130_fd_sc_hd__o2bb2ai_4 _14988_ (.A1_N(_10519_),
    .A2_N(_10530_),
    .B1(_10552_),
    .B2(_09390_),
    .Y(_10607_));
 sky130_fd_sc_hd__nand3_4 _14989_ (.A(_10574_),
    .B(_10530_),
    .C(_10519_),
    .Y(_10618_));
 sky130_fd_sc_hd__a22oi_1 _14990_ (.A1(_06804_),
    .A2(_06826_),
    .B1(_10585_),
    .B2(_10596_),
    .Y(_10629_));
 sky130_fd_sc_hd__nand3_1 _14991_ (.A(_10607_),
    .B(_10618_),
    .C(_06837_),
    .Y(_10640_));
 sky130_fd_sc_hd__a31oi_4 _14992_ (.A1(_10607_),
    .A2(_10618_),
    .A3(_06837_),
    .B1(_10486_),
    .Y(_10651_));
 sky130_fd_sc_hd__o21ai_1 _14993_ (.A1(_08568_),
    .A2(_09511_),
    .B1(_09631_),
    .Y(_10662_));
 sky130_fd_sc_hd__a22oi_1 _14994_ (.A1(_08579_),
    .A2(_09522_),
    .B1(_09489_),
    .B2(net385),
    .Y(_10673_));
 sky130_fd_sc_hd__a21oi_1 _14995_ (.A1(_09533_),
    .A2(_09631_),
    .B1(_09642_),
    .Y(_10684_));
 sky130_fd_sc_hd__o21ai_1 _14996_ (.A1(net385),
    .A2(_09489_),
    .B1(_10662_),
    .Y(_10695_));
 sky130_fd_sc_hd__a31o_1 _14997_ (.A1(_10607_),
    .A2(_10618_),
    .A3(_06837_),
    .B1(_05862_),
    .X(_10706_));
 sky130_fd_sc_hd__a311oi_4 _14998_ (.A1(_10607_),
    .A2(_10618_),
    .A3(_06837_),
    .B1(_10486_),
    .C1(_05862_),
    .Y(_10717_));
 sky130_fd_sc_hd__o211ai_1 _14999_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_10497_),
    .C1(_10640_),
    .Y(_10728_));
 sky130_fd_sc_hd__a2bb2oi_1 _15000_ (.A1_N(_05763_),
    .A2_N(_05785_),
    .B1(_10497_),
    .B2(_10640_),
    .Y(_10739_));
 sky130_fd_sc_hd__o22ai_2 _15001_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_10486_),
    .B2(_10629_),
    .Y(_10750_));
 sky130_fd_sc_hd__o211ai_1 _15002_ (.A1(_09642_),
    .A2(_10673_),
    .B1(_10728_),
    .C1(_10750_),
    .Y(_10761_));
 sky130_fd_sc_hd__o21ai_1 _15003_ (.A1(_10717_),
    .A2(_10739_),
    .B1(_10684_),
    .Y(_10772_));
 sky130_fd_sc_hd__nand3_2 _15004_ (.A(_10772_),
    .B(_07713_),
    .C(_10761_),
    .Y(_10783_));
 sky130_fd_sc_hd__o21ai_4 _15005_ (.A1(_07713_),
    .A2(_10651_),
    .B1(_10783_),
    .Y(_10794_));
 sky130_fd_sc_hd__a31oi_4 _15006_ (.A1(_05250_),
    .A2(_09587_),
    .A3(_09609_),
    .B1(_08645_),
    .Y(_10805_));
 sky130_fd_sc_hd__nand2_1 _15007_ (.A(_09675_),
    .B(_08634_),
    .Y(_10816_));
 sky130_fd_sc_hd__a2bb2oi_1 _15008_ (.A1_N(net398),
    .A2_N(net397),
    .B1(_09697_),
    .B2(_10816_),
    .Y(_10827_));
 sky130_fd_sc_hd__o22ai_4 _15009_ (.A1(net398),
    .A2(net397),
    .B1(_09686_),
    .B2(_10805_),
    .Y(_10838_));
 sky130_fd_sc_hd__o211ai_4 _15010_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_09697_),
    .C1(_10816_),
    .Y(_10849_));
 sky130_fd_sc_hd__a31oi_2 _15011_ (.A1(_10838_),
    .A2(_10849_),
    .A3(_08721_),
    .B1(_10794_),
    .Y(_10860_));
 sky130_fd_sc_hd__a31o_1 _15012_ (.A1(_10838_),
    .A2(_10849_),
    .A3(_08721_),
    .B1(_10794_),
    .X(_10871_));
 sky130_fd_sc_hd__nand4_2 _15013_ (.A(_10838_),
    .B(_08721_),
    .C(_10794_),
    .D(_10849_),
    .Y(_10882_));
 sky130_fd_sc_hd__o221ai_2 _15014_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_07713_),
    .B2(_10651_),
    .C1(_10783_),
    .Y(_10893_));
 sky130_fd_sc_hd__o21ai_2 _15015_ (.A1(net398),
    .A2(net397),
    .B1(_10794_),
    .Y(_10904_));
 sky130_fd_sc_hd__a41oi_4 _15016_ (.A1(_08721_),
    .A2(_10794_),
    .A3(_10838_),
    .A4(_10849_),
    .B1(_10860_),
    .Y(_10915_));
 sky130_fd_sc_hd__a21oi_1 _15017_ (.A1(_10871_),
    .A2(_10882_),
    .B1(net403),
    .Y(_10926_));
 sky130_fd_sc_hd__a21o_1 _15018_ (.A1(_10871_),
    .A2(_10882_),
    .B1(net403),
    .X(_10937_));
 sky130_fd_sc_hd__nand3_4 _15019_ (.A(_10871_),
    .B(_10882_),
    .C(net403),
    .Y(_10948_));
 sky130_fd_sc_hd__a21o_1 _15020_ (.A1(_10937_),
    .A2(_10948_),
    .B1(_09862_),
    .X(_10959_));
 sky130_fd_sc_hd__o211ai_1 _15021_ (.A1(_09730_),
    .A2(_03289_),
    .B1(_10948_),
    .C1(_10937_),
    .Y(_10969_));
 sky130_fd_sc_hd__nand3_1 _15022_ (.A(_10959_),
    .B(_10969_),
    .C(_09829_),
    .Y(_10980_));
 sky130_fd_sc_hd__o31a_1 _15023_ (.A1(net350),
    .A2(net349),
    .A3(_10915_),
    .B1(_10980_),
    .X(_10991_));
 sky130_fd_sc_hd__o311a_4 _15024_ (.A1(net350),
    .A2(net349),
    .A3(_10915_),
    .B1(net1),
    .C1(_10980_),
    .X(_11002_));
 sky130_fd_sc_hd__o211ai_1 _15025_ (.A1(_09829_),
    .A2(_10915_),
    .B1(net1),
    .C1(_10980_),
    .Y(_11013_));
 sky130_fd_sc_hd__nor2_1 _15026_ (.A(net1),
    .B(_10991_),
    .Y(_11024_));
 sky130_fd_sc_hd__o41a_1 _15027_ (.A1(net60),
    .A2(net61),
    .A3(net62),
    .A4(_07680_),
    .B1(net409),
    .X(_11035_));
 sky130_fd_sc_hd__and2b_4 _15028_ (.A_N(_11035_),
    .B(net63),
    .X(_11046_));
 sky130_fd_sc_hd__and2b_4 _15029_ (.A_N(net63),
    .B(_11035_),
    .X(_11057_));
 sky130_fd_sc_hd__or2_4 _15030_ (.A(net347),
    .B(net346),
    .X(_11068_));
 sky130_fd_sc_hd__nor2_8 _15031_ (.A(net347),
    .B(net346),
    .Y(_11079_));
 sky130_fd_sc_hd__o21ai_1 _15032_ (.A1(_11002_),
    .A2(_11024_),
    .B1(_11068_),
    .Y(_11090_));
 sky130_fd_sc_hd__o31a_2 _15033_ (.A1(_10991_),
    .A2(net347),
    .A3(net346),
    .B1(_11090_),
    .X(_11101_));
 sky130_fd_sc_hd__a21oi_1 _15034_ (.A1(_05119_),
    .A2(_09894_),
    .B1(_11101_),
    .Y(_11112_));
 sky130_fd_sc_hd__and3_1 _15035_ (.A(_05119_),
    .B(_09894_),
    .C(_11101_),
    .X(_11123_));
 sky130_fd_sc_hd__nor2_1 _15036_ (.A(_11112_),
    .B(_11123_),
    .Y(net127));
 sky130_fd_sc_hd__o22a_1 _15037_ (.A1(_04832_),
    .A2(_04942_),
    .B1(_09894_),
    .B2(_11101_),
    .X(_11144_));
 sky130_fd_sc_hd__o211a_1 _15038_ (.A1(_09379_),
    .A2(_09390_),
    .B1(_09423_),
    .C1(_10519_),
    .X(_11155_));
 sky130_fd_sc_hd__o211ai_1 _15039_ (.A1(_09379_),
    .A2(_09390_),
    .B1(_09423_),
    .C1(_10519_),
    .Y(_11166_));
 sky130_fd_sc_hd__o21a_1 _15040_ (.A1(_10508_),
    .A2(_10574_),
    .B1(_10530_),
    .X(_11177_));
 sky130_fd_sc_hd__o21ai_4 _15041_ (.A1(_10508_),
    .A2(_10574_),
    .B1(_10530_),
    .Y(_11188_));
 sky130_fd_sc_hd__o21ai_2 _15042_ (.A1(net31),
    .A2(_09916_),
    .B1(net410),
    .Y(_11199_));
 sky130_fd_sc_hd__o311a_4 _15043_ (.A1(net30),
    .A2(net31),
    .A3(_08808_),
    .B1(_04172_),
    .C1(net410),
    .X(_11210_));
 sky130_fd_sc_hd__or2_2 _15044_ (.A(net32),
    .B(_11199_),
    .X(_11221_));
 sky130_fd_sc_hd__and2_4 _15045_ (.A(_11199_),
    .B(net32),
    .X(_11232_));
 sky130_fd_sc_hd__nand2_2 _15046_ (.A(_11199_),
    .B(net32),
    .Y(_11243_));
 sky130_fd_sc_hd__o311a_4 _15047_ (.A1(net30),
    .A2(net31),
    .A3(_08808_),
    .B1(net32),
    .C1(net410),
    .X(_11254_));
 sky130_fd_sc_hd__o211ai_4 _15048_ (.A1(net31),
    .A2(_09916_),
    .B1(net32),
    .C1(net410),
    .Y(_11265_));
 sky130_fd_sc_hd__and2_4 _15049_ (.A(_04172_),
    .B(_11199_),
    .X(_11276_));
 sky130_fd_sc_hd__clkinv_4 _15050_ (.A(_11276_),
    .Y(_11287_));
 sky130_fd_sc_hd__nor2_8 _15051_ (.A(_11210_),
    .B(_11232_),
    .Y(_11298_));
 sky130_fd_sc_hd__nor2_8 _15052_ (.A(_11254_),
    .B(_11276_),
    .Y(_11309_));
 sky130_fd_sc_hd__o21a_2 _15053_ (.A1(_11210_),
    .A2(_11232_),
    .B1(net33),
    .X(_11320_));
 sky130_fd_sc_hd__o32a_2 _15054_ (.A1(_03178_),
    .A2(_11254_),
    .A3(_11276_),
    .B1(net408),
    .B2(_05152_),
    .X(_11331_));
 sky130_fd_sc_hd__a31o_1 _15055_ (.A1(_11287_),
    .A2(net33),
    .A3(_11265_),
    .B1(net404),
    .X(_11342_));
 sky130_fd_sc_hd__and3_1 _15056_ (.A(net330),
    .B(net33),
    .C(net348),
    .X(_11353_));
 sky130_fd_sc_hd__or4_1 _15057_ (.A(_03178_),
    .B(_09971_),
    .C(_09993_),
    .D(net331),
    .X(_11364_));
 sky130_fd_sc_hd__o32a_1 _15058_ (.A1(_03178_),
    .A2(_11254_),
    .A3(_11276_),
    .B1(_09971_),
    .B2(net363),
    .X(_11375_));
 sky130_fd_sc_hd__a31o_1 _15059_ (.A1(_11287_),
    .A2(net33),
    .A3(_11265_),
    .B1(net348),
    .X(_11386_));
 sky130_fd_sc_hd__o21ai_1 _15060_ (.A1(_10036_),
    .A2(net331),
    .B1(_11386_),
    .Y(_11397_));
 sky130_fd_sc_hd__o2111ai_2 _15061_ (.A1(_07077_),
    .A2(_07888_),
    .B1(_07942_),
    .C1(_07121_),
    .D1(_07143_),
    .Y(_11408_));
 sky130_fd_sc_hd__nor2_2 _15062_ (.A(_08951_),
    .B(_11408_),
    .Y(_11419_));
 sky130_fd_sc_hd__and3_4 _15063_ (.A(_07187_),
    .B(_10113_),
    .C(_11419_),
    .X(_11430_));
 sky130_fd_sc_hd__o2111ai_4 _15064_ (.A1(_10015_),
    .A2(_08929_),
    .B1(_07187_),
    .C1(_10080_),
    .D1(_11419_),
    .Y(_11441_));
 sky130_fd_sc_hd__o2bb2a_1 _15065_ (.A1_N(_10080_),
    .A2_N(_11419_),
    .B1(_08929_),
    .B2(_10015_),
    .X(_11452_));
 sky130_fd_sc_hd__a32o_1 _15066_ (.A1(net33),
    .A2(_08918_),
    .A3(net348),
    .B1(_11419_),
    .B2(_10080_),
    .X(_11463_));
 sky130_fd_sc_hd__a21oi_4 _15067_ (.A1(_10069_),
    .A2(_10113_),
    .B1(_11463_),
    .Y(_11473_));
 sky130_fd_sc_hd__o21ai_2 _15068_ (.A1(_10124_),
    .A2(_10058_),
    .B1(_11452_),
    .Y(_11484_));
 sky130_fd_sc_hd__a31o_1 _15069_ (.A1(_07187_),
    .A2(_10113_),
    .A3(_11419_),
    .B1(_11473_),
    .X(_11495_));
 sky130_fd_sc_hd__inv_2 _15070_ (.A(_11495_),
    .Y(_11506_));
 sky130_fd_sc_hd__nor3_1 _15071_ (.A(_11397_),
    .B(_11430_),
    .C(_11473_),
    .Y(_11517_));
 sky130_fd_sc_hd__o2111ai_4 _15072_ (.A1(_10036_),
    .A2(net331),
    .B1(_11386_),
    .C1(_11441_),
    .D1(_11484_),
    .Y(_11528_));
 sky130_fd_sc_hd__o22a_1 _15073_ (.A1(_11353_),
    .A2(_11375_),
    .B1(_11430_),
    .B2(_11473_),
    .X(_11539_));
 sky130_fd_sc_hd__o22ai_4 _15074_ (.A1(_11353_),
    .A2(_11375_),
    .B1(_11430_),
    .B2(_11473_),
    .Y(_11550_));
 sky130_fd_sc_hd__nand2_2 _15075_ (.A(_11528_),
    .B(_11550_),
    .Y(_11561_));
 sky130_fd_sc_hd__a21oi_4 _15076_ (.A1(_11528_),
    .A2(_11550_),
    .B1(_05185_),
    .Y(_11572_));
 sky130_fd_sc_hd__o21bai_1 _15077_ (.A1(_11517_),
    .A2(_11539_),
    .B1_N(_05185_),
    .Y(_11583_));
 sky130_fd_sc_hd__a21oi_4 _15078_ (.A1(_11561_),
    .A2(net404),
    .B1(_11331_),
    .Y(_11594_));
 sky130_fd_sc_hd__a31oi_4 _15079_ (.A1(_09094_),
    .A2(_10245_),
    .A3(_10267_),
    .B1(_10256_),
    .Y(_11605_));
 sky130_fd_sc_hd__a31o_2 _15080_ (.A1(_09094_),
    .A2(_10245_),
    .A3(_10267_),
    .B1(_10256_),
    .X(_11616_));
 sky130_fd_sc_hd__or3_4 _15081_ (.A(_08863_),
    .B(net366),
    .C(_11331_),
    .X(_11627_));
 sky130_fd_sc_hd__a21oi_2 _15082_ (.A1(_11561_),
    .A2(net404),
    .B1(_11627_),
    .Y(_11638_));
 sky130_fd_sc_hd__a21o_1 _15083_ (.A1(_11561_),
    .A2(net404),
    .B1(_11627_),
    .X(_11649_));
 sky130_fd_sc_hd__a2bb2oi_2 _15084_ (.A1_N(_08863_),
    .A2_N(net366),
    .B1(_11342_),
    .B2(_11583_),
    .Y(_11660_));
 sky130_fd_sc_hd__o22ai_4 _15085_ (.A1(_08863_),
    .A2(net366),
    .B1(_11331_),
    .B2(_11572_),
    .Y(_11671_));
 sky130_fd_sc_hd__o21ai_1 _15086_ (.A1(_11572_),
    .A2(_11627_),
    .B1(_11671_),
    .Y(_11682_));
 sky130_fd_sc_hd__o211a_1 _15087_ (.A1(_11627_),
    .A2(_11572_),
    .B1(_11616_),
    .C1(_11671_),
    .X(_11693_));
 sky130_fd_sc_hd__o211ai_4 _15088_ (.A1(_11627_),
    .A2(_11572_),
    .B1(_11616_),
    .C1(_11671_),
    .Y(_11704_));
 sky130_fd_sc_hd__a21oi_1 _15089_ (.A1(_11649_),
    .A2(_11671_),
    .B1(_11616_),
    .Y(_11715_));
 sky130_fd_sc_hd__o21bai_1 _15090_ (.A1(_11638_),
    .A2(_11660_),
    .B1_N(_11616_),
    .Y(_11726_));
 sky130_fd_sc_hd__o22ai_4 _15091_ (.A1(net402),
    .A2(net399),
    .B1(_11693_),
    .B2(_11715_),
    .Y(_11737_));
 sky130_fd_sc_hd__or4_2 _15092_ (.A(net402),
    .B(net399),
    .C(_11331_),
    .D(_11572_),
    .X(_11748_));
 sky130_fd_sc_hd__a22oi_4 _15093_ (.A1(_05359_),
    .A2(_05381_),
    .B1(_11682_),
    .B2(_11605_),
    .Y(_11759_));
 sky130_fd_sc_hd__o211ai_2 _15094_ (.A1(net402),
    .A2(net399),
    .B1(_11704_),
    .C1(_11726_),
    .Y(_11770_));
 sky130_fd_sc_hd__a22o_2 _15095_ (.A1(_05392_),
    .A2(_11594_),
    .B1(_11759_),
    .B2(_11704_),
    .X(_11781_));
 sky130_fd_sc_hd__a22oi_4 _15096_ (.A1(_05392_),
    .A2(_11594_),
    .B1(_11759_),
    .B2(_11704_),
    .Y(_11792_));
 sky130_fd_sc_hd__o221a_2 _15097_ (.A1(_05654_),
    .A2(_05665_),
    .B1(_11594_),
    .B2(net388),
    .C1(_11737_),
    .X(_11803_));
 sky130_fd_sc_hd__or3_1 _15098_ (.A(net384),
    .B(net383),
    .C(_11792_),
    .X(_11814_));
 sky130_fd_sc_hd__a2bb2oi_1 _15099_ (.A1_N(net389),
    .A2_N(net370),
    .B1(_11748_),
    .B2(_11770_),
    .Y(_11825_));
 sky130_fd_sc_hd__o211ai_4 _15100_ (.A1(_11594_),
    .A2(net388),
    .B1(_07899_),
    .C1(_11737_),
    .Y(_11836_));
 sky130_fd_sc_hd__o211ai_4 _15101_ (.A1(net369),
    .A2(_07866_),
    .B1(_11748_),
    .C1(_11770_),
    .Y(_11847_));
 sky130_fd_sc_hd__nor2_2 _15102_ (.A(_10366_),
    .B(_10388_),
    .Y(_11858_));
 sky130_fd_sc_hd__o21ai_4 _15103_ (.A1(_10355_),
    .A2(_10399_),
    .B1(_10377_),
    .Y(_11869_));
 sky130_fd_sc_hd__a21oi_2 _15104_ (.A1(_11836_),
    .A2(_11847_),
    .B1(_11869_),
    .Y(_11880_));
 sky130_fd_sc_hd__o2bb2ai_4 _15105_ (.A1_N(_11836_),
    .A2_N(_11847_),
    .B1(_11858_),
    .B2(_10355_),
    .Y(_11891_));
 sky130_fd_sc_hd__nand3_2 _15106_ (.A(_11836_),
    .B(_11847_),
    .C(_11869_),
    .Y(_11902_));
 sky130_fd_sc_hd__a31oi_2 _15107_ (.A1(_11836_),
    .A2(_11847_),
    .A3(_11869_),
    .B1(_05731_),
    .Y(_11913_));
 sky130_fd_sc_hd__a31o_1 _15108_ (.A1(_11836_),
    .A2(_11847_),
    .A3(_11869_),
    .B1(_05731_),
    .X(_11924_));
 sky130_fd_sc_hd__nand3_1 _15109_ (.A(_11891_),
    .B(_11902_),
    .C(net360),
    .Y(_11935_));
 sky130_fd_sc_hd__a22oi_4 _15110_ (.A1(_05731_),
    .A2(_11781_),
    .B1(_11913_),
    .B2(_11891_),
    .Y(_11946_));
 sky130_fd_sc_hd__o22ai_4 _15111_ (.A1(net360),
    .A2(_11792_),
    .B1(_11880_),
    .B2(_11924_),
    .Y(_11956_));
 sky130_fd_sc_hd__a31o_1 _15112_ (.A1(_11891_),
    .A2(_11902_),
    .A3(net360),
    .B1(_07044_),
    .X(_11967_));
 sky130_fd_sc_hd__a311oi_4 _15113_ (.A1(_11891_),
    .A2(_11902_),
    .A3(net360),
    .B1(_07044_),
    .C1(_11803_),
    .Y(_11978_));
 sky130_fd_sc_hd__o221ai_4 _15114_ (.A1(net360),
    .A2(_11792_),
    .B1(_11880_),
    .B2(_11924_),
    .C1(_07033_),
    .Y(_11989_));
 sky130_fd_sc_hd__a2bb2oi_1 _15115_ (.A1_N(_06945_),
    .A2_N(net377),
    .B1(_11814_),
    .B2(_11935_),
    .Y(_12000_));
 sky130_fd_sc_hd__o21ai_2 _15116_ (.A1(_06945_),
    .A2(net377),
    .B1(_11956_),
    .Y(_12011_));
 sky130_fd_sc_hd__nand3_2 _15117_ (.A(_12011_),
    .B(_11177_),
    .C(_11989_),
    .Y(_12022_));
 sky130_fd_sc_hd__o22ai_4 _15118_ (.A1(_10541_),
    .A2(_11155_),
    .B1(_11978_),
    .B2(_12000_),
    .Y(_12033_));
 sky130_fd_sc_hd__and3_1 _15119_ (.A(_06804_),
    .B(_06826_),
    .C(_11956_),
    .X(_12044_));
 sky130_fd_sc_hd__or3_2 _15120_ (.A(net379),
    .B(net378),
    .C(_11946_),
    .X(_12055_));
 sky130_fd_sc_hd__nand3_4 _15121_ (.A(_12033_),
    .B(_06837_),
    .C(_12022_),
    .Y(_12066_));
 sky130_fd_sc_hd__o21ai_1 _15122_ (.A1(_06837_),
    .A2(_11946_),
    .B1(_12066_),
    .Y(_12077_));
 sky130_fd_sc_hd__a31oi_2 _15123_ (.A1(_12033_),
    .A2(_06837_),
    .A3(_12022_),
    .B1(_12044_),
    .Y(_12088_));
 sky130_fd_sc_hd__a21oi_2 _15124_ (.A1(_12055_),
    .A2(_12066_),
    .B1(_07713_),
    .Y(_12099_));
 sky130_fd_sc_hd__or3_2 _15125_ (.A(net372),
    .B(net371),
    .C(_12088_),
    .X(_12110_));
 sky130_fd_sc_hd__a2bb2oi_2 _15126_ (.A1_N(net393),
    .A2_N(net382),
    .B1(_12055_),
    .B2(_12066_),
    .Y(_12121_));
 sky130_fd_sc_hd__a22o_1 _15127_ (.A1(_06256_),
    .A2(_06278_),
    .B1(_12055_),
    .B2(_12066_),
    .X(_12132_));
 sky130_fd_sc_hd__o221a_1 _15128_ (.A1(net380),
    .A2(net391),
    .B1(_06837_),
    .B2(_11946_),
    .C1(_12066_),
    .X(_12143_));
 sky130_fd_sc_hd__o221ai_4 _15129_ (.A1(net380),
    .A2(net391),
    .B1(_06837_),
    .B2(_11946_),
    .C1(_12066_),
    .Y(_12154_));
 sky130_fd_sc_hd__o221a_1 _15130_ (.A1(_09620_),
    .A2(_09544_),
    .B1(_05851_),
    .B2(_10651_),
    .C1(_09653_),
    .X(_12165_));
 sky130_fd_sc_hd__a2bb2oi_2 _15131_ (.A1_N(_10486_),
    .A2_N(_10706_),
    .B1(_10684_),
    .B2(_10750_),
    .Y(_12176_));
 sky130_fd_sc_hd__o22ai_2 _15132_ (.A1(_10486_),
    .A2(_10706_),
    .B1(_10739_),
    .B2(_10695_),
    .Y(_12187_));
 sky130_fd_sc_hd__o21ai_2 _15133_ (.A1(_12121_),
    .A2(_12143_),
    .B1(_12187_),
    .Y(_12198_));
 sky130_fd_sc_hd__nand3_2 _15134_ (.A(_12132_),
    .B(_12154_),
    .C(_12176_),
    .Y(_12209_));
 sky130_fd_sc_hd__nand3_2 _15135_ (.A(_12198_),
    .B(_12209_),
    .C(_07713_),
    .Y(_12220_));
 sky130_fd_sc_hd__a31oi_4 _15136_ (.A1(_12198_),
    .A2(_12209_),
    .A3(_07713_),
    .B1(_12099_),
    .Y(_12231_));
 sky130_fd_sc_hd__a31o_1 _15137_ (.A1(_12198_),
    .A2(_12209_),
    .A3(_07713_),
    .B1(_12099_),
    .X(_12242_));
 sky130_fd_sc_hd__o21ai_2 _15138_ (.A1(_09686_),
    .A2(_10805_),
    .B1(_10893_),
    .Y(_12253_));
 sky130_fd_sc_hd__nand2_1 _15139_ (.A(_12253_),
    .B(_10904_),
    .Y(_12264_));
 sky130_fd_sc_hd__o21ai_1 _15140_ (.A1(_10794_),
    .A2(_10827_),
    .B1(_10849_),
    .Y(_12275_));
 sky130_fd_sc_hd__o211ai_4 _15141_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_10904_),
    .C1(_12253_),
    .Y(_12286_));
 sky130_fd_sc_hd__o211ai_2 _15142_ (.A1(_10794_),
    .A2(_10827_),
    .B1(_10849_),
    .C1(_05862_),
    .Y(_12297_));
 sky130_fd_sc_hd__a21oi_2 _15143_ (.A1(_12264_),
    .A2(_05862_),
    .B1(_08732_),
    .Y(_12308_));
 sky130_fd_sc_hd__and4_2 _15144_ (.A(_12297_),
    .B(_08721_),
    .C(_12286_),
    .D(_12231_),
    .X(_12319_));
 sky130_fd_sc_hd__a31oi_4 _15145_ (.A1(_12297_),
    .A2(_08721_),
    .A3(_12286_),
    .B1(_12231_),
    .Y(_12330_));
 sky130_fd_sc_hd__a2bb2oi_1 _15146_ (.A1_N(_05763_),
    .A2_N(_05785_),
    .B1(_12110_),
    .B2(_12220_),
    .Y(_12341_));
 sky130_fd_sc_hd__a22o_1 _15147_ (.A1(_05774_),
    .A2(_05796_),
    .B1(_12110_),
    .B2(_12220_),
    .X(_12352_));
 sky130_fd_sc_hd__nand3_1 _15148_ (.A(_12220_),
    .B(_05851_),
    .C(_12110_),
    .Y(_12363_));
 sky130_fd_sc_hd__nand2_1 _15149_ (.A(_12363_),
    .B(_12264_),
    .Y(_12374_));
 sky130_fd_sc_hd__a41oi_4 _15150_ (.A1(_12220_),
    .A2(_12308_),
    .A3(_12286_),
    .A4(_12110_),
    .B1(_12330_),
    .Y(_12385_));
 sky130_fd_sc_hd__a41o_1 _15151_ (.A1(_12220_),
    .A2(_12308_),
    .A3(_12286_),
    .A4(_12110_),
    .B1(_12330_),
    .X(_12396_));
 sky130_fd_sc_hd__o21ai_4 _15152_ (.A1(_03289_),
    .A2(_09730_),
    .B1(_10948_),
    .Y(_12407_));
 sky130_fd_sc_hd__o21ai_1 _15153_ (.A1(net403),
    .A2(_10915_),
    .B1(_12407_),
    .Y(_12417_));
 sky130_fd_sc_hd__and3_1 _15154_ (.A(_05556_),
    .B(_10937_),
    .C(_12407_),
    .X(_12428_));
 sky130_fd_sc_hd__o211ai_4 _15155_ (.A1(net398),
    .A2(net397),
    .B1(_10937_),
    .C1(_12407_),
    .Y(_12439_));
 sky130_fd_sc_hd__o221ai_4 _15156_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_09862_),
    .B2(_10926_),
    .C1(_10948_),
    .Y(_12450_));
 sky130_fd_sc_hd__nand3_1 _15157_ (.A(_12450_),
    .B(_09829_),
    .C(_12439_),
    .Y(_12461_));
 sky130_fd_sc_hd__a31o_1 _15158_ (.A1(_12450_),
    .A2(_09829_),
    .A3(_12439_),
    .B1(_12396_),
    .X(_12472_));
 sky130_fd_sc_hd__nand4_4 _15159_ (.A(_12396_),
    .B(_12439_),
    .C(_12450_),
    .D(_09829_),
    .Y(_12483_));
 sky130_fd_sc_hd__nand4_4 _15160_ (.A(_12450_),
    .B(_12385_),
    .C(_09829_),
    .D(_12439_),
    .Y(_12494_));
 sky130_fd_sc_hd__o21ai_4 _15161_ (.A1(_12319_),
    .A2(_12330_),
    .B1(_12461_),
    .Y(_12505_));
 sky130_fd_sc_hd__o21ai_1 _15162_ (.A1(_12319_),
    .A2(_12330_),
    .B1(_05556_),
    .Y(_12516_));
 sky130_fd_sc_hd__nand2_1 _15163_ (.A(_12472_),
    .B(_12483_),
    .Y(_12527_));
 sky130_fd_sc_hd__a21oi_2 _15164_ (.A1(_12494_),
    .A2(_12505_),
    .B1(_05250_),
    .Y(_12538_));
 sky130_fd_sc_hd__nand4_2 _15165_ (.A(_05207_),
    .B(_05229_),
    .C(_12472_),
    .D(_12483_),
    .Y(_12549_));
 sky130_fd_sc_hd__nand3_4 _15166_ (.A(_05250_),
    .B(_12494_),
    .C(_12505_),
    .Y(_12560_));
 sky130_fd_sc_hd__a21oi_1 _15167_ (.A1(_12549_),
    .A2(_12560_),
    .B1(_11002_),
    .Y(_12571_));
 sky130_fd_sc_hd__a31oi_2 _15168_ (.A1(_05250_),
    .A2(_12494_),
    .A3(_12505_),
    .B1(_11013_),
    .Y(_12582_));
 sky130_fd_sc_hd__nand2_1 _15169_ (.A(_12560_),
    .B(_11002_),
    .Y(_12593_));
 sky130_fd_sc_hd__a31o_1 _15170_ (.A1(_12549_),
    .A2(_12560_),
    .A3(_11002_),
    .B1(_11079_),
    .X(_12604_));
 sky130_fd_sc_hd__o22ai_2 _15171_ (.A1(_11068_),
    .A2(_12527_),
    .B1(_12571_),
    .B2(_12604_),
    .Y(_12615_));
 sky130_fd_sc_hd__and2_1 _15172_ (.A(net1),
    .B(_12615_),
    .X(_12626_));
 sky130_fd_sc_hd__nand2_2 _15173_ (.A(net1),
    .B(_12615_),
    .Y(_12637_));
 sky130_fd_sc_hd__o221a_1 _15174_ (.A1(_11068_),
    .A2(_12527_),
    .B1(_12571_),
    .B2(_12604_),
    .C1(_03289_),
    .X(_12648_));
 sky130_fd_sc_hd__or3_4 _15175_ (.A(net62),
    .B(net63),
    .C(_09752_),
    .X(_12659_));
 sky130_fd_sc_hd__a21boi_4 _15176_ (.A1(_12659_),
    .A2(net409),
    .B1_N(net64),
    .Y(_12670_));
 sky130_fd_sc_hd__and3b_4 _15177_ (.A_N(net64),
    .B(_12659_),
    .C(net409),
    .X(_12681_));
 sky130_fd_sc_hd__or2_4 _15178_ (.A(net328),
    .B(_12681_),
    .X(_12692_));
 sky130_fd_sc_hd__nor2_8 _15179_ (.A(net328),
    .B(_12681_),
    .Y(_12703_));
 sky130_fd_sc_hd__o21ai_1 _15180_ (.A1(_12626_),
    .A2(_12648_),
    .B1(_12692_),
    .Y(_12714_));
 sky130_fd_sc_hd__o31a_1 _15181_ (.A1(_12615_),
    .A2(net328),
    .A3(_12681_),
    .B1(_12714_),
    .X(_12725_));
 sky130_fd_sc_hd__xor2_1 _15182_ (.A(_11144_),
    .B(_12725_),
    .X(net128));
 sky130_fd_sc_hd__nor3_1 _15183_ (.A(_09894_),
    .B(_11101_),
    .C(_12725_),
    .Y(_12746_));
 sky130_fd_sc_hd__o31a_1 _15184_ (.A1(_09894_),
    .A2(_11101_),
    .A3(_12725_),
    .B1(_05119_),
    .X(_12757_));
 sky130_fd_sc_hd__a21oi_1 _15185_ (.A1(_12077_),
    .A2(_06343_),
    .B1(_12176_),
    .Y(_12768_));
 sky130_fd_sc_hd__o22ai_4 _15186_ (.A1(_10717_),
    .A2(_12165_),
    .B1(_06332_),
    .B2(_12088_),
    .Y(_12779_));
 sky130_fd_sc_hd__a31oi_2 _15187_ (.A1(_06332_),
    .A2(_12055_),
    .A3(_12066_),
    .B1(_12187_),
    .Y(_12790_));
 sky130_fd_sc_hd__a21oi_1 _15188_ (.A1(_12154_),
    .A2(_12176_),
    .B1(_12121_),
    .Y(_12801_));
 sky130_fd_sc_hd__nor2_1 _15189_ (.A(net31),
    .B(net32),
    .Y(_12812_));
 sky130_fd_sc_hd__or2_2 _15190_ (.A(net31),
    .B(net32),
    .X(_12823_));
 sky130_fd_sc_hd__and4b_2 _15191_ (.A_N(_07789_),
    .B(_12812_),
    .C(_03952_),
    .D(_04062_),
    .X(_12834_));
 sky130_fd_sc_hd__o311a_4 _15192_ (.A1(_12823_),
    .A2(net30),
    .A3(_08808_),
    .B1(_04282_),
    .C1(net410),
    .X(_12845_));
 sky130_fd_sc_hd__o21a_4 _15193_ (.A1(_03399_),
    .A2(_12834_),
    .B1(net2),
    .X(_12856_));
 sky130_fd_sc_hd__o21a_4 _15194_ (.A1(_03399_),
    .A2(_12834_),
    .B1(_04282_),
    .X(_12867_));
 sky130_fd_sc_hd__o311a_4 _15195_ (.A1(_12823_),
    .A2(net30),
    .A3(_08808_),
    .B1(net2),
    .C1(net410),
    .X(_12877_));
 sky130_fd_sc_hd__nor2_8 _15196_ (.A(net361),
    .B(net345),
    .Y(_12888_));
 sky130_fd_sc_hd__nor2_8 _15197_ (.A(_12867_),
    .B(_12877_),
    .Y(_12899_));
 sky130_fd_sc_hd__or3_4 _15198_ (.A(_12877_),
    .B(_03178_),
    .C(_12867_),
    .X(_12910_));
 sky130_fd_sc_hd__and3_1 _15199_ (.A(net325),
    .B(net33),
    .C(net330),
    .X(_12921_));
 sky130_fd_sc_hd__or4_2 _15200_ (.A(_03178_),
    .B(_11254_),
    .C(_11276_),
    .D(_12888_),
    .X(_12932_));
 sky130_fd_sc_hd__o32a_1 _15201_ (.A1(_12877_),
    .A2(_03178_),
    .A3(_12867_),
    .B1(_11254_),
    .B2(_11276_),
    .X(_12943_));
 sky130_fd_sc_hd__or4_1 _15202_ (.A(_03178_),
    .B(_12867_),
    .C(_12877_),
    .D(net330),
    .X(_12954_));
 sky130_fd_sc_hd__a22o_1 _15203_ (.A1(_11221_),
    .A2(_11243_),
    .B1(net326),
    .B2(net33),
    .X(_12965_));
 sky130_fd_sc_hd__a21oi_2 _15204_ (.A1(_11320_),
    .A2(net325),
    .B1(_12943_),
    .Y(_12976_));
 sky130_fd_sc_hd__a21o_1 _15205_ (.A1(_11320_),
    .A2(net325),
    .B1(_12943_),
    .X(_12987_));
 sky130_fd_sc_hd__o22ai_4 _15206_ (.A1(_10036_),
    .A2(net331),
    .B1(_11430_),
    .B2(_11473_),
    .Y(_12998_));
 sky130_fd_sc_hd__o21a_1 _15207_ (.A1(net348),
    .A2(_11320_),
    .B1(_11441_),
    .X(_13009_));
 sky130_fd_sc_hd__a21boi_1 _15208_ (.A1(_10146_),
    .A2(_11452_),
    .B1_N(_13009_),
    .Y(_13020_));
 sky130_fd_sc_hd__nand2_1 _15209_ (.A(_11484_),
    .B(_13009_),
    .Y(_13031_));
 sky130_fd_sc_hd__nor3_1 _15210_ (.A(_11353_),
    .B(_12976_),
    .C(_13020_),
    .Y(_13042_));
 sky130_fd_sc_hd__o211ai_2 _15211_ (.A1(_10036_),
    .A2(net331),
    .B1(_12987_),
    .C1(_13031_),
    .Y(_13053_));
 sky130_fd_sc_hd__a22oi_2 _15212_ (.A1(_12954_),
    .A2(_12965_),
    .B1(_13031_),
    .B2(_11364_),
    .Y(_13064_));
 sky130_fd_sc_hd__o211ai_4 _15213_ (.A1(net348),
    .A2(_11320_),
    .B1(_12976_),
    .C1(_12998_),
    .Y(_13075_));
 sky130_fd_sc_hd__nand3_2 _15214_ (.A(_13075_),
    .B(net404),
    .C(_13053_),
    .Y(_13086_));
 sky130_fd_sc_hd__o32a_1 _15215_ (.A1(_12877_),
    .A2(_03178_),
    .A3(_12867_),
    .B1(net408),
    .B2(_05152_),
    .X(_13097_));
 sky130_fd_sc_hd__a21oi_2 _15216_ (.A1(_13053_),
    .A2(_13075_),
    .B1(_05185_),
    .Y(_13108_));
 sky130_fd_sc_hd__o21ai_1 _15217_ (.A1(_13042_),
    .A2(_13064_),
    .B1(net404),
    .Y(_13119_));
 sky130_fd_sc_hd__o21ai_4 _15218_ (.A1(net404),
    .A2(_12910_),
    .B1(_13086_),
    .Y(_13130_));
 sky130_fd_sc_hd__a211o_2 _15219_ (.A1(_05185_),
    .A2(_12910_),
    .B1(net388),
    .C1(_13108_),
    .X(_13141_));
 sky130_fd_sc_hd__inv_2 _15220_ (.A(_13141_),
    .Y(_13152_));
 sky130_fd_sc_hd__a21oi_4 _15221_ (.A1(_11616_),
    .A2(_11671_),
    .B1(_11638_),
    .Y(_13163_));
 sky130_fd_sc_hd__o21ai_2 _15222_ (.A1(_11605_),
    .A2(_11660_),
    .B1(_11649_),
    .Y(_13174_));
 sky130_fd_sc_hd__o221ai_4 _15223_ (.A1(_09971_),
    .A2(net363),
    .B1(_12910_),
    .B2(net404),
    .C1(_13086_),
    .Y(_13185_));
 sky130_fd_sc_hd__a21oi_1 _15224_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_13097_),
    .Y(_13196_));
 sky130_fd_sc_hd__or3_2 _15225_ (.A(_09971_),
    .B(net363),
    .C(_13097_),
    .X(_13207_));
 sky130_fd_sc_hd__nand2_2 _15226_ (.A(_13119_),
    .B(_13196_),
    .Y(_13218_));
 sky130_fd_sc_hd__o21a_2 _15227_ (.A1(_13207_),
    .A2(_13108_),
    .B1(_13185_),
    .X(_13229_));
 sky130_fd_sc_hd__o21ai_4 _15228_ (.A1(_13207_),
    .A2(_13108_),
    .B1(_13185_),
    .Y(_13240_));
 sky130_fd_sc_hd__o211ai_2 _15229_ (.A1(_11572_),
    .A2(_11627_),
    .B1(_11704_),
    .C1(_13240_),
    .Y(_13251_));
 sky130_fd_sc_hd__nand2_2 _15230_ (.A(_13174_),
    .B(_13229_),
    .Y(_13262_));
 sky130_fd_sc_hd__nand2_1 _15231_ (.A(_13163_),
    .B(_13229_),
    .Y(_13273_));
 sky130_fd_sc_hd__a22oi_4 _15232_ (.A1(_05359_),
    .A2(_05381_),
    .B1(_13163_),
    .B2(_13240_),
    .Y(_13284_));
 sky130_fd_sc_hd__o211a_1 _15233_ (.A1(_13240_),
    .A2(_13163_),
    .B1(net388),
    .C1(_13251_),
    .X(_13295_));
 sky130_fd_sc_hd__o211ai_2 _15234_ (.A1(_13240_),
    .A2(_13163_),
    .B1(net388),
    .C1(_13251_),
    .Y(_13306_));
 sky130_fd_sc_hd__a22oi_4 _15235_ (.A1(_05392_),
    .A2(_13130_),
    .B1(_13284_),
    .B2(_13262_),
    .Y(_13317_));
 sky130_fd_sc_hd__a22o_1 _15236_ (.A1(_05392_),
    .A2(_13130_),
    .B1(_13284_),
    .B2(_13262_),
    .X(_13328_));
 sky130_fd_sc_hd__o22ai_4 _15237_ (.A1(_10355_),
    .A2(_11858_),
    .B1(_07888_),
    .B2(_11792_),
    .Y(_13339_));
 sky130_fd_sc_hd__nand2_1 _15238_ (.A(_11847_),
    .B(_11869_),
    .Y(_13349_));
 sky130_fd_sc_hd__a21oi_2 _15239_ (.A1(_11847_),
    .A2(_11869_),
    .B1(_11825_),
    .Y(_13360_));
 sky130_fd_sc_hd__and3_2 _15240_ (.A(_05687_),
    .B(_05709_),
    .C(_13328_),
    .X(_13371_));
 sky130_fd_sc_hd__or3_2 _15241_ (.A(net384),
    .B(net383),
    .C(_13317_),
    .X(_13382_));
 sky130_fd_sc_hd__a21oi_1 _15242_ (.A1(_13284_),
    .A2(_13262_),
    .B1(_08918_),
    .Y(_13393_));
 sky130_fd_sc_hd__o311a_2 _15243_ (.A1(net388),
    .A2(_13097_),
    .A3(_13108_),
    .B1(_08907_),
    .C1(_13306_),
    .X(_13404_));
 sky130_fd_sc_hd__nand3_2 _15244_ (.A(_13306_),
    .B(_08907_),
    .C(_13141_),
    .Y(_13415_));
 sky130_fd_sc_hd__a21oi_1 _15245_ (.A1(_13141_),
    .A2(_13306_),
    .B1(_08907_),
    .Y(_13426_));
 sky130_fd_sc_hd__o22ai_4 _15246_ (.A1(_08819_),
    .A2(net367),
    .B1(_13152_),
    .B2(_13295_),
    .Y(_13437_));
 sky130_fd_sc_hd__o2111ai_4 _15247_ (.A1(_11781_),
    .A2(_07899_),
    .B1(_13415_),
    .C1(_13339_),
    .D1(_13437_),
    .Y(_13448_));
 sky130_fd_sc_hd__o2bb2ai_4 _15248_ (.A1_N(_11847_),
    .A2_N(_13339_),
    .B1(_13404_),
    .B2(_13426_),
    .Y(_13459_));
 sky130_fd_sc_hd__o211ai_4 _15249_ (.A1(net384),
    .A2(net383),
    .B1(_13448_),
    .C1(_13459_),
    .Y(_13470_));
 sky130_fd_sc_hd__a31oi_4 _15250_ (.A1(_13448_),
    .A2(_13459_),
    .A3(net360),
    .B1(_13371_),
    .Y(_13481_));
 sky130_fd_sc_hd__a31o_1 _15251_ (.A1(_13448_),
    .A2(_13459_),
    .A3(net360),
    .B1(_13371_),
    .X(_13492_));
 sky130_fd_sc_hd__and3_2 _15252_ (.A(_06804_),
    .B(_06826_),
    .C(_13492_),
    .X(_13503_));
 sky130_fd_sc_hd__or3_4 _15253_ (.A(net379),
    .B(net378),
    .C(_13481_),
    .X(_13514_));
 sky130_fd_sc_hd__a22oi_2 _15254_ (.A1(_10530_),
    .A2(_11166_),
    .B1(_11956_),
    .B2(_07044_),
    .Y(_13525_));
 sky130_fd_sc_hd__o21ai_4 _15255_ (.A1(_07033_),
    .A2(_11946_),
    .B1(_11188_),
    .Y(_13536_));
 sky130_fd_sc_hd__o21ai_1 _15256_ (.A1(_11188_),
    .A2(_11978_),
    .B1(_12011_),
    .Y(_13547_));
 sky130_fd_sc_hd__a311oi_4 _15257_ (.A1(_13448_),
    .A2(_13459_),
    .A3(net360),
    .B1(_07899_),
    .C1(_13371_),
    .Y(_13558_));
 sky130_fd_sc_hd__nand3_4 _15258_ (.A(_13470_),
    .B(_07888_),
    .C(_13382_),
    .Y(_13569_));
 sky130_fd_sc_hd__a22oi_4 _15259_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_13382_),
    .B2(_13470_),
    .Y(_13580_));
 sky130_fd_sc_hd__o211ai_4 _15260_ (.A1(_11967_),
    .A2(_11803_),
    .B1(_13569_),
    .C1(_13536_),
    .Y(_13591_));
 sky130_fd_sc_hd__o311ai_4 _15261_ (.A1(net369),
    .A2(_07866_),
    .A3(_13481_),
    .B1(_13569_),
    .C1(_13547_),
    .Y(_13602_));
 sky130_fd_sc_hd__o22ai_4 _15262_ (.A1(_11978_),
    .A2(_13525_),
    .B1(_13558_),
    .B2(_13580_),
    .Y(_13613_));
 sky130_fd_sc_hd__o211a_1 _15263_ (.A1(_13580_),
    .A2(_13591_),
    .B1(_06837_),
    .C1(_13613_),
    .X(_13624_));
 sky130_fd_sc_hd__o211ai_4 _15264_ (.A1(_13580_),
    .A2(_13591_),
    .B1(_06837_),
    .C1(_13613_),
    .Y(_13635_));
 sky130_fd_sc_hd__a31oi_4 _15265_ (.A1(_13602_),
    .A2(_13613_),
    .A3(_06837_),
    .B1(_13503_),
    .Y(_13646_));
 sky130_fd_sc_hd__a31o_1 _15266_ (.A1(_13602_),
    .A2(_13613_),
    .A3(_06837_),
    .B1(_13503_),
    .X(_13657_));
 sky130_fd_sc_hd__a311oi_4 _15267_ (.A1(_13602_),
    .A2(_13613_),
    .A3(_06837_),
    .B1(_07044_),
    .C1(_13503_),
    .Y(_13668_));
 sky130_fd_sc_hd__nand3_4 _15268_ (.A(_13635_),
    .B(_07033_),
    .C(_13514_),
    .Y(_13679_));
 sky130_fd_sc_hd__a2bb2oi_4 _15269_ (.A1_N(_06945_),
    .A2_N(net377),
    .B1(_13514_),
    .B2(_13635_),
    .Y(_13690_));
 sky130_fd_sc_hd__o22ai_4 _15270_ (.A1(_06945_),
    .A2(net377),
    .B1(_13503_),
    .B2(_13624_),
    .Y(_13701_));
 sky130_fd_sc_hd__o211ai_4 _15271_ (.A1(_12121_),
    .A2(_12790_),
    .B1(_13679_),
    .C1(_13701_),
    .Y(_13712_));
 sky130_fd_sc_hd__o22ai_4 _15272_ (.A1(_12143_),
    .A2(_12768_),
    .B1(_13668_),
    .B2(_13690_),
    .Y(_13723_));
 sky130_fd_sc_hd__a21oi_4 _15273_ (.A1(_13514_),
    .A2(_13635_),
    .B1(_07713_),
    .Y(_13734_));
 sky130_fd_sc_hd__or3_2 _15274_ (.A(net372),
    .B(net371),
    .C(_13646_),
    .X(_13745_));
 sky130_fd_sc_hd__o211a_1 _15275_ (.A1(net372),
    .A2(net371),
    .B1(_13712_),
    .C1(_13723_),
    .X(_13756_));
 sky130_fd_sc_hd__o211ai_4 _15276_ (.A1(net372),
    .A2(net371),
    .B1(_13712_),
    .C1(_13723_),
    .Y(_13767_));
 sky130_fd_sc_hd__a31o_1 _15277_ (.A1(_13712_),
    .A2(_13723_),
    .A3(_07713_),
    .B1(_13734_),
    .X(_13778_));
 sky130_fd_sc_hd__a31oi_4 _15278_ (.A1(_13712_),
    .A2(_13723_),
    .A3(_07713_),
    .B1(_13734_),
    .Y(_13788_));
 sky130_fd_sc_hd__and3_1 _15279_ (.A(_13778_),
    .B(_08711_),
    .C(_08689_),
    .X(_13799_));
 sky130_fd_sc_hd__a2bb2oi_4 _15280_ (.A1_N(net393),
    .A2_N(net382),
    .B1(_13745_),
    .B2(_13767_),
    .Y(_13810_));
 sky130_fd_sc_hd__o22ai_2 _15281_ (.A1(net392),
    .A2(net382),
    .B1(_13734_),
    .B2(_13756_),
    .Y(_13821_));
 sky130_fd_sc_hd__o221a_1 _15282_ (.A1(net380),
    .A2(net391),
    .B1(_07713_),
    .B2(_13646_),
    .C1(_13767_),
    .X(_13832_));
 sky130_fd_sc_hd__nand3_2 _15283_ (.A(_13767_),
    .B(_06332_),
    .C(_13745_),
    .Y(_13843_));
 sky130_fd_sc_hd__o21ai_1 _15284_ (.A1(_05851_),
    .A2(_12231_),
    .B1(_12275_),
    .Y(_13854_));
 sky130_fd_sc_hd__a21oi_2 _15285_ (.A1(_12363_),
    .A2(_12264_),
    .B1(_12341_),
    .Y(_13865_));
 sky130_fd_sc_hd__o2bb2ai_2 _15286_ (.A1_N(_12352_),
    .A2_N(_12374_),
    .B1(_13810_),
    .B2(_13832_),
    .Y(_13876_));
 sky130_fd_sc_hd__nand3_2 _15287_ (.A(_13821_),
    .B(_13843_),
    .C(_13865_),
    .Y(_13887_));
 sky130_fd_sc_hd__o21ai_2 _15288_ (.A1(_13810_),
    .A2(_13832_),
    .B1(_13865_),
    .Y(_13898_));
 sky130_fd_sc_hd__a22oi_1 _15289_ (.A1(_13788_),
    .A2(_06332_),
    .B1(_12352_),
    .B2(_12374_),
    .Y(_13909_));
 sky130_fd_sc_hd__o211ai_4 _15290_ (.A1(_05862_),
    .A2(_12242_),
    .B1(_13843_),
    .C1(_13854_),
    .Y(_13920_));
 sky130_fd_sc_hd__o221a_1 _15291_ (.A1(net353),
    .A2(net352),
    .B1(_13810_),
    .B2(_13920_),
    .C1(_13898_),
    .X(_13931_));
 sky130_fd_sc_hd__o221ai_4 _15292_ (.A1(net353),
    .A2(net352),
    .B1(_13810_),
    .B2(_13920_),
    .C1(_13898_),
    .Y(_13942_));
 sky130_fd_sc_hd__nand3_2 _15293_ (.A(_13876_),
    .B(_13887_),
    .C(_08721_),
    .Y(_13953_));
 sky130_fd_sc_hd__o311a_1 _15294_ (.A1(net372),
    .A2(net371),
    .A3(_13646_),
    .B1(_13767_),
    .C1(_08732_),
    .X(_13964_));
 sky130_fd_sc_hd__or4_1 _15295_ (.A(net353),
    .B(net352),
    .C(_13734_),
    .D(_13756_),
    .X(_13975_));
 sky130_fd_sc_hd__o31a_1 _15296_ (.A1(_08721_),
    .A2(_13734_),
    .A3(_13756_),
    .B1(_13953_),
    .X(_13986_));
 sky130_fd_sc_hd__a2bb2oi_2 _15297_ (.A1_N(_12319_),
    .A2_N(_12330_),
    .B1(net385),
    .B2(_12417_),
    .Y(_13997_));
 sky130_fd_sc_hd__o221ai_4 _15298_ (.A1(net403),
    .A2(_10915_),
    .B1(_12319_),
    .B2(_12330_),
    .C1(_12407_),
    .Y(_14008_));
 sky130_fd_sc_hd__a21boi_1 _15299_ (.A1(_12396_),
    .A2(_12450_),
    .B1_N(_12439_),
    .Y(_14019_));
 sky130_fd_sc_hd__o211ai_4 _15300_ (.A1(net385),
    .A2(_12385_),
    .B1(_12439_),
    .C1(_14008_),
    .Y(_14030_));
 sky130_fd_sc_hd__and4_1 _15301_ (.A(_12439_),
    .B(_12516_),
    .C(_14008_),
    .D(_05851_),
    .X(_14041_));
 sky130_fd_sc_hd__o2111ai_2 _15302_ (.A1(net385),
    .A2(_12417_),
    .B1(_12516_),
    .C1(_05851_),
    .D1(_14008_),
    .Y(_14052_));
 sky130_fd_sc_hd__o22ai_2 _15303_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_12428_),
    .B2(_13997_),
    .Y(_14063_));
 sky130_fd_sc_hd__a31oi_2 _15304_ (.A1(_14063_),
    .A2(_09829_),
    .A3(_14052_),
    .B1(_13986_),
    .Y(_14074_));
 sky130_fd_sc_hd__o2111a_1 _15305_ (.A1(_13799_),
    .A2(_13931_),
    .B1(_09829_),
    .C1(_14052_),
    .D1(_14063_),
    .X(_14085_));
 sky130_fd_sc_hd__o221a_1 _15306_ (.A1(_09763_),
    .A2(_09774_),
    .B1(_13778_),
    .B2(_08721_),
    .C1(_13953_),
    .X(_14096_));
 sky130_fd_sc_hd__a311o_1 _15307_ (.A1(_13876_),
    .A2(_13887_),
    .A3(_08721_),
    .B1(_13964_),
    .C1(_09829_),
    .X(_14107_));
 sky130_fd_sc_hd__a311oi_4 _15308_ (.A1(_13876_),
    .A2(_13887_),
    .A3(_08721_),
    .B1(_13964_),
    .C1(_05851_),
    .Y(_14118_));
 sky130_fd_sc_hd__o211ai_2 _15309_ (.A1(_08721_),
    .A2(_13778_),
    .B1(_13953_),
    .C1(_05862_),
    .Y(_14129_));
 sky130_fd_sc_hd__a21oi_1 _15310_ (.A1(_13953_),
    .A2(_13975_),
    .B1(_05862_),
    .Y(_14140_));
 sky130_fd_sc_hd__o221ai_4 _15311_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_08721_),
    .B2(_13788_),
    .C1(_13942_),
    .Y(_14151_));
 sky130_fd_sc_hd__o211ai_4 _15312_ (.A1(_12428_),
    .A2(_13997_),
    .B1(_14129_),
    .C1(_14151_),
    .Y(_14162_));
 sky130_fd_sc_hd__o21ai_2 _15313_ (.A1(_14118_),
    .A2(_14140_),
    .B1(_14019_),
    .Y(_14173_));
 sky130_fd_sc_hd__nand3_1 _15314_ (.A(_14173_),
    .B(_09829_),
    .C(_14162_),
    .Y(_14184_));
 sky130_fd_sc_hd__a31o_2 _15315_ (.A1(_14173_),
    .A2(_09829_),
    .A3(_14162_),
    .B1(_14096_),
    .X(_14195_));
 sky130_fd_sc_hd__a31oi_4 _15316_ (.A1(_14173_),
    .A2(_09829_),
    .A3(_14162_),
    .B1(_14096_),
    .Y(_14206_));
 sky130_fd_sc_hd__a32oi_4 _15317_ (.A1(net403),
    .A2(_12472_),
    .A3(_12483_),
    .B1(_12560_),
    .B2(_11002_),
    .Y(_14216_));
 sky130_fd_sc_hd__a221oi_4 _15318_ (.A1(_05512_),
    .A2(_05534_),
    .B1(_12560_),
    .B2(_11002_),
    .C1(_12538_),
    .Y(_14227_));
 sky130_fd_sc_hd__nand3_4 _15319_ (.A(_12593_),
    .B(net385),
    .C(_12549_),
    .Y(_14238_));
 sky130_fd_sc_hd__o22ai_4 _15320_ (.A1(net398),
    .A2(net397),
    .B1(_12538_),
    .B2(_12582_),
    .Y(_14249_));
 sky130_fd_sc_hd__o211ai_2 _15321_ (.A1(net347),
    .A2(net346),
    .B1(_14238_),
    .C1(_14249_),
    .Y(_14260_));
 sky130_fd_sc_hd__o2111a_2 _15322_ (.A1(net347),
    .A2(net346),
    .B1(_14238_),
    .C1(_14249_),
    .D1(_14195_),
    .X(_14271_));
 sky130_fd_sc_hd__o2111ai_4 _15323_ (.A1(net347),
    .A2(net346),
    .B1(_14238_),
    .C1(_14249_),
    .D1(_14195_),
    .Y(_14282_));
 sky130_fd_sc_hd__a31oi_4 _15324_ (.A1(_14249_),
    .A2(_11068_),
    .A3(_14238_),
    .B1(_14195_),
    .Y(_14293_));
 sky130_fd_sc_hd__o21ai_1 _15325_ (.A1(_14074_),
    .A2(_14085_),
    .B1(_14260_),
    .Y(_14304_));
 sky130_fd_sc_hd__a211oi_2 _15326_ (.A1(_05458_),
    .A2(_05480_),
    .B1(_14074_),
    .C1(_14085_),
    .Y(_14315_));
 sky130_fd_sc_hd__a31o_1 _15327_ (.A1(_14107_),
    .A2(_14184_),
    .A3(_14260_),
    .B1(_14271_),
    .X(_14326_));
 sky130_fd_sc_hd__a311o_2 _15328_ (.A1(_14107_),
    .A2(_14184_),
    .A3(_14260_),
    .B1(_05250_),
    .C1(_14271_),
    .X(_14337_));
 sky130_fd_sc_hd__a21oi_4 _15329_ (.A1(_14282_),
    .A2(_14304_),
    .B1(net403),
    .Y(_14348_));
 sky130_fd_sc_hd__o21ai_1 _15330_ (.A1(_14271_),
    .A2(_14293_),
    .B1(_05250_),
    .Y(_14359_));
 sky130_fd_sc_hd__a21oi_1 _15331_ (.A1(_14337_),
    .A2(_14359_),
    .B1(_12626_),
    .Y(_14370_));
 sky130_fd_sc_hd__nand2_1 _15332_ (.A(_14359_),
    .B(_12626_),
    .Y(_14381_));
 sky130_fd_sc_hd__a31o_1 _15333_ (.A1(_14337_),
    .A2(_14359_),
    .A3(_12626_),
    .B1(_12703_),
    .X(_14392_));
 sky130_fd_sc_hd__o22ai_2 _15334_ (.A1(_12692_),
    .A2(_14326_),
    .B1(_14370_),
    .B2(_14392_),
    .Y(_14403_));
 sky130_fd_sc_hd__and2_2 _15335_ (.A(net1),
    .B(_14403_),
    .X(_14414_));
 sky130_fd_sc_hd__nand2_2 _15336_ (.A(net1),
    .B(_14403_),
    .Y(_14425_));
 sky130_fd_sc_hd__o221a_1 _15337_ (.A1(_12692_),
    .A2(_14326_),
    .B1(_14370_),
    .B2(_14392_),
    .C1(_03289_),
    .X(_14436_));
 sky130_fd_sc_hd__or4_4 _15338_ (.A(net62),
    .B(net63),
    .C(net64),
    .D(_09752_),
    .X(_14447_));
 sky130_fd_sc_hd__and3_4 _15339_ (.A(_14447_),
    .B(net34),
    .C(net409),
    .X(_14458_));
 sky130_fd_sc_hd__a21oi_4 _15340_ (.A1(_14447_),
    .A2(net409),
    .B1(net34),
    .Y(_00000_));
 sky130_fd_sc_hd__and3b_4 _15341_ (.A_N(net34),
    .B(_14447_),
    .C(net409),
    .X(_00011_));
 sky130_fd_sc_hd__inv_2 _15342_ (.A(_00011_),
    .Y(_00022_));
 sky130_fd_sc_hd__a21boi_4 _15343_ (.A1(_14447_),
    .A2(net409),
    .B1_N(net34),
    .Y(_00033_));
 sky130_fd_sc_hd__inv_2 _15344_ (.A(net321),
    .Y(_00044_));
 sky130_fd_sc_hd__nor2_4 _15345_ (.A(_14458_),
    .B(_00000_),
    .Y(_00055_));
 sky130_fd_sc_hd__nor2_8 _15346_ (.A(net324),
    .B(net322),
    .Y(_00066_));
 sky130_fd_sc_hd__o21ai_1 _15347_ (.A1(_14458_),
    .A2(_00000_),
    .B1(_14403_),
    .Y(_00077_));
 sky130_fd_sc_hd__o31a_1 _15348_ (.A1(_00066_),
    .A2(_14436_),
    .A3(_14414_),
    .B1(_00077_),
    .X(_00088_));
 sky130_fd_sc_hd__xnor2_1 _15349_ (.A(_12757_),
    .B(_00088_),
    .Y(net66));
 sky130_fd_sc_hd__a2bb2o_1 _15350_ (.A1_N(_04832_),
    .A2_N(_04942_),
    .B1(_12746_),
    .B2(_00088_),
    .X(_00109_));
 sky130_fd_sc_hd__a2bb2oi_1 _15351_ (.A1_N(_07888_),
    .A2_N(_13481_),
    .B1(_13536_),
    .B2(_11989_),
    .Y(_00120_));
 sky130_fd_sc_hd__o221ai_4 _15352_ (.A1(_11978_),
    .A2(_11188_),
    .B1(_07888_),
    .B2(_13481_),
    .C1(_12011_),
    .Y(_00131_));
 sky130_fd_sc_hd__a31oi_4 _15353_ (.A1(_11989_),
    .A2(_13536_),
    .A3(_13569_),
    .B1(_13580_),
    .Y(_00142_));
 sky130_fd_sc_hd__and3_1 _15354_ (.A(_09905_),
    .B(_12812_),
    .C(_04282_),
    .X(_00152_));
 sky130_fd_sc_hd__or4_4 _15355_ (.A(net30),
    .B(_12823_),
    .C(net2),
    .D(_08808_),
    .X(_00163_));
 sky130_fd_sc_hd__o311a_4 _15356_ (.A1(_12823_),
    .A2(net2),
    .A3(_09916_),
    .B1(_04392_),
    .C1(net410),
    .X(_00174_));
 sky130_fd_sc_hd__a311o_4 _15357_ (.A1(_09905_),
    .A2(_12812_),
    .A3(_04282_),
    .B1(net3),
    .C1(_03399_),
    .X(_00185_));
 sky130_fd_sc_hd__a21oi_4 _15358_ (.A1(_00163_),
    .A2(net410),
    .B1(_04392_),
    .Y(_00196_));
 sky130_fd_sc_hd__a21o_4 _15359_ (.A1(_00163_),
    .A2(net410),
    .B1(_04392_),
    .X(_00207_));
 sky130_fd_sc_hd__a21oi_4 _15360_ (.A1(_00163_),
    .A2(net410),
    .B1(net3),
    .Y(_00218_));
 sky130_fd_sc_hd__o311a_4 _15361_ (.A1(_12823_),
    .A2(net2),
    .A3(_09916_),
    .B1(net3),
    .C1(net410),
    .X(_00229_));
 sky130_fd_sc_hd__nor2_8 _15362_ (.A(_00174_),
    .B(net344),
    .Y(_00240_));
 sky130_fd_sc_hd__nor2_8 _15363_ (.A(_00218_),
    .B(_00229_),
    .Y(_00251_));
 sky130_fd_sc_hd__o21a_1 _15364_ (.A1(_00174_),
    .A2(_00196_),
    .B1(net33),
    .X(_00262_));
 sky130_fd_sc_hd__or3_4 _15365_ (.A(_03178_),
    .B(_00218_),
    .C(_00229_),
    .X(_00273_));
 sky130_fd_sc_hd__a31oi_2 _15366_ (.A1(_11386_),
    .A2(_12998_),
    .A3(_12976_),
    .B1(_12921_),
    .Y(_00284_));
 sky130_fd_sc_hd__or3_1 _15367_ (.A(_12845_),
    .B(_12856_),
    .C(_00262_),
    .X(_00295_));
 sky130_fd_sc_hd__o21ai_4 _15368_ (.A1(_12910_),
    .A2(net320),
    .B1(_00295_),
    .Y(_00306_));
 sky130_fd_sc_hd__a21oi_4 _15369_ (.A1(_12932_),
    .A2(_13075_),
    .B1(_00306_),
    .Y(_00317_));
 sky130_fd_sc_hd__o21bai_2 _15370_ (.A1(_12921_),
    .A2(_13064_),
    .B1_N(_00306_),
    .Y(_00328_));
 sky130_fd_sc_hd__o211ai_4 _15371_ (.A1(_12910_),
    .A2(net331),
    .B1(_00306_),
    .C1(_13075_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_2 _15372_ (.A(_00339_),
    .B(_05174_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand3_1 _15373_ (.A(_00328_),
    .B(_00339_),
    .C(_05174_),
    .Y(_00361_));
 sky130_fd_sc_hd__o221a_1 _15374_ (.A1(net408),
    .A2(_05152_),
    .B1(_00174_),
    .B2(_00196_),
    .C1(net33),
    .X(_00372_));
 sky130_fd_sc_hd__or4_2 _15375_ (.A(_03178_),
    .B(_05174_),
    .C(_00218_),
    .D(_00229_),
    .X(_00383_));
 sky130_fd_sc_hd__o22ai_4 _15376_ (.A1(net404),
    .A2(_00273_),
    .B1(_00317_),
    .B2(_00350_),
    .Y(_00394_));
 sky130_fd_sc_hd__o32a_2 _15377_ (.A1(_03178_),
    .A2(net404),
    .A3(net320),
    .B1(_00317_),
    .B2(_00350_),
    .X(_00405_));
 sky130_fd_sc_hd__or3_2 _15378_ (.A(net402),
    .B(net400),
    .C(_00405_),
    .X(_00416_));
 sky130_fd_sc_hd__a311oi_4 _15379_ (.A1(_00328_),
    .A2(_00339_),
    .A3(_05174_),
    .B1(_00372_),
    .C1(net330),
    .Y(_00427_));
 sky130_fd_sc_hd__o221ai_4 _15380_ (.A1(net404),
    .A2(_00273_),
    .B1(_00317_),
    .B2(_00350_),
    .C1(net331),
    .Y(_00438_));
 sky130_fd_sc_hd__a21oi_4 _15381_ (.A1(_00361_),
    .A2(_00383_),
    .B1(net331),
    .Y(_00449_));
 sky130_fd_sc_hd__o21ai_2 _15382_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_00394_),
    .Y(_00460_));
 sky130_fd_sc_hd__nor2_2 _15383_ (.A(_00427_),
    .B(_00449_),
    .Y(_00471_));
 sky130_fd_sc_hd__o211ai_4 _15384_ (.A1(_11605_),
    .A2(_11660_),
    .B1(_13218_),
    .C1(_11649_),
    .Y(_00482_));
 sky130_fd_sc_hd__o2111a_1 _15385_ (.A1(net348),
    .A2(_13130_),
    .B1(_00438_),
    .C1(_00460_),
    .D1(_00482_),
    .X(_00493_));
 sky130_fd_sc_hd__o2111ai_4 _15386_ (.A1(net348),
    .A2(_13130_),
    .B1(_00438_),
    .C1(_00460_),
    .D1(_00482_),
    .Y(_00504_));
 sky130_fd_sc_hd__o211a_1 _15387_ (.A1(_00427_),
    .A2(_00449_),
    .B1(_13218_),
    .C1(_13262_),
    .X(_00515_));
 sky130_fd_sc_hd__o211ai_2 _15388_ (.A1(_00427_),
    .A2(_00449_),
    .B1(_13218_),
    .C1(_13262_),
    .Y(_00525_));
 sky130_fd_sc_hd__o211ai_4 _15389_ (.A1(net402),
    .A2(net399),
    .B1(_00504_),
    .C1(_00525_),
    .Y(_00536_));
 sky130_fd_sc_hd__o311a_1 _15390_ (.A1(_03178_),
    .A2(_05174_),
    .A3(net320),
    .B1(_05392_),
    .C1(_00361_),
    .X(_00547_));
 sky130_fd_sc_hd__a21oi_1 _15391_ (.A1(_00504_),
    .A2(_00525_),
    .B1(_05392_),
    .Y(_00558_));
 sky130_fd_sc_hd__o22ai_2 _15392_ (.A1(net402),
    .A2(net399),
    .B1(_00493_),
    .B2(_00515_),
    .Y(_00569_));
 sky130_fd_sc_hd__o31a_1 _15393_ (.A1(net402),
    .A2(net400),
    .A3(_00405_),
    .B1(_00536_),
    .X(_00580_));
 sky130_fd_sc_hd__o21ai_2 _15394_ (.A1(net388),
    .A2(_00405_),
    .B1(_00536_),
    .Y(_00591_));
 sky130_fd_sc_hd__o311a_1 _15395_ (.A1(net402),
    .A2(_00405_),
    .A3(net400),
    .B1(_05731_),
    .C1(_00536_),
    .X(_00602_));
 sky130_fd_sc_hd__a2bb2oi_4 _15396_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_00416_),
    .B2(_00536_),
    .Y(_00613_));
 sky130_fd_sc_hd__o221ai_4 _15397_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_00394_),
    .B2(net388),
    .C1(_00569_),
    .Y(_00624_));
 sky130_fd_sc_hd__o211a_1 _15398_ (.A1(net388),
    .A2(_00405_),
    .B1(_10015_),
    .C1(_00536_),
    .X(_00635_));
 sky130_fd_sc_hd__nand3_4 _15399_ (.A(_00536_),
    .B(_10015_),
    .C(_00416_),
    .Y(_00646_));
 sky130_fd_sc_hd__o221ai_4 _15400_ (.A1(_11792_),
    .A2(_07888_),
    .B1(_08907_),
    .B2(_13317_),
    .C1(_13349_),
    .Y(_00657_));
 sky130_fd_sc_hd__a22oi_4 _15401_ (.A1(_13393_),
    .A2(_13141_),
    .B1(_13360_),
    .B2(_13437_),
    .Y(_00668_));
 sky130_fd_sc_hd__o21ai_1 _15402_ (.A1(_08918_),
    .A2(_13328_),
    .B1(_00657_),
    .Y(_00679_));
 sky130_fd_sc_hd__o2111ai_4 _15403_ (.A1(_13360_),
    .A2(_13404_),
    .B1(_13437_),
    .C1(_00624_),
    .D1(_00646_),
    .Y(_00690_));
 sky130_fd_sc_hd__o21ai_2 _15404_ (.A1(_00613_),
    .A2(_00635_),
    .B1(_00668_),
    .Y(_00701_));
 sky130_fd_sc_hd__o211ai_2 _15405_ (.A1(net384),
    .A2(net383),
    .B1(_00690_),
    .C1(_00701_),
    .Y(_00712_));
 sky130_fd_sc_hd__o221a_2 _15406_ (.A1(_05654_),
    .A2(_05665_),
    .B1(_00394_),
    .B2(net388),
    .C1(_00569_),
    .X(_00723_));
 sky130_fd_sc_hd__o21ai_4 _15407_ (.A1(_00613_),
    .A2(_00635_),
    .B1(_00679_),
    .Y(_00734_));
 sky130_fd_sc_hd__o211ai_4 _15408_ (.A1(_08918_),
    .A2(_13328_),
    .B1(_00646_),
    .C1(_00657_),
    .Y(_00745_));
 sky130_fd_sc_hd__o211ai_4 _15409_ (.A1(net348),
    .A2(_00591_),
    .B1(_00624_),
    .C1(_00668_),
    .Y(_00756_));
 sky130_fd_sc_hd__o211ai_1 _15410_ (.A1(_00613_),
    .A2(_00745_),
    .B1(_05720_),
    .C1(_00734_),
    .Y(_00767_));
 sky130_fd_sc_hd__a31oi_4 _15411_ (.A1(_00734_),
    .A2(_00756_),
    .A3(_05720_),
    .B1(_00723_),
    .Y(_00778_));
 sky130_fd_sc_hd__a311oi_4 _15412_ (.A1(_00734_),
    .A2(_00756_),
    .A3(_05720_),
    .B1(_08918_),
    .C1(_00723_),
    .Y(_00789_));
 sky130_fd_sc_hd__o211ai_2 _15413_ (.A1(_05720_),
    .A2(_00580_),
    .B1(_08907_),
    .C1(_00767_),
    .Y(_00800_));
 sky130_fd_sc_hd__a311oi_4 _15414_ (.A1(_00690_),
    .A2(_00701_),
    .A3(net360),
    .B1(_08907_),
    .C1(_00602_),
    .Y(_00811_));
 sky130_fd_sc_hd__o211ai_2 _15415_ (.A1(_00591_),
    .A2(net360),
    .B1(_08918_),
    .C1(_00712_),
    .Y(_00822_));
 sky130_fd_sc_hd__o2111ai_4 _15416_ (.A1(_07899_),
    .A2(_13492_),
    .B1(_00131_),
    .C1(_00800_),
    .D1(_00822_),
    .Y(_00833_));
 sky130_fd_sc_hd__o22ai_4 _15417_ (.A1(_13558_),
    .A2(_00120_),
    .B1(_00789_),
    .B2(_00811_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand3_4 _15418_ (.A(_00844_),
    .B(_06837_),
    .C(_00833_),
    .Y(_00855_));
 sky130_fd_sc_hd__o211a_1 _15419_ (.A1(_00591_),
    .A2(net360),
    .B1(_06848_),
    .C1(_00712_),
    .X(_00866_));
 sky130_fd_sc_hd__a311o_4 _15420_ (.A1(_00690_),
    .A2(_00701_),
    .A3(net360),
    .B1(_06837_),
    .C1(_00602_),
    .X(_00877_));
 sky130_fd_sc_hd__a31o_1 _15421_ (.A1(_00844_),
    .A2(_06837_),
    .A3(_00833_),
    .B1(_00866_),
    .X(_00888_));
 sky130_fd_sc_hd__a31oi_4 _15422_ (.A1(_00844_),
    .A2(_06837_),
    .A3(_00833_),
    .B1(_00866_),
    .Y(_00899_));
 sky130_fd_sc_hd__o311a_1 _15423_ (.A1(net379),
    .A2(_00778_),
    .A3(net378),
    .B1(_07724_),
    .C1(_00855_),
    .X(_00910_));
 sky130_fd_sc_hd__a22oi_4 _15424_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_00855_),
    .B2(_00877_),
    .Y(_00920_));
 sky130_fd_sc_hd__a22o_2 _15425_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_00855_),
    .B2(_00877_),
    .X(_00931_));
 sky130_fd_sc_hd__o221a_1 _15426_ (.A1(net369),
    .A2(_07866_),
    .B1(_00778_),
    .B2(_06837_),
    .C1(_00855_),
    .X(_00942_));
 sky130_fd_sc_hd__nand3_4 _15427_ (.A(_00855_),
    .B(_00877_),
    .C(_07888_),
    .Y(_00953_));
 sky130_fd_sc_hd__o21ai_2 _15428_ (.A1(_07033_),
    .A2(_13646_),
    .B1(_12801_),
    .Y(_00964_));
 sky130_fd_sc_hd__o211ai_1 _15429_ (.A1(_12077_),
    .A2(_06343_),
    .B1(_13679_),
    .C1(_12779_),
    .Y(_00975_));
 sky130_fd_sc_hd__o21bai_1 _15430_ (.A1(_13668_),
    .A2(_12801_),
    .B1_N(_13690_),
    .Y(_00986_));
 sky130_fd_sc_hd__a31oi_4 _15431_ (.A1(_12154_),
    .A2(_12779_),
    .A3(_13679_),
    .B1(_13690_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand3_1 _15432_ (.A(_00931_),
    .B(_00953_),
    .C(_00997_),
    .Y(_01008_));
 sky130_fd_sc_hd__o21ai_1 _15433_ (.A1(_00920_),
    .A2(_00942_),
    .B1(_00986_),
    .Y(_01019_));
 sky130_fd_sc_hd__o21ai_4 _15434_ (.A1(_00920_),
    .A2(_00942_),
    .B1(_00997_),
    .Y(_01030_));
 sky130_fd_sc_hd__a22oi_2 _15435_ (.A1(_00899_),
    .A2(_07888_),
    .B1(_13701_),
    .B2(_00975_),
    .Y(_01041_));
 sky130_fd_sc_hd__o211ai_4 _15436_ (.A1(_07044_),
    .A2(_13657_),
    .B1(_00953_),
    .C1(_00964_),
    .Y(_01052_));
 sky130_fd_sc_hd__nand3_2 _15437_ (.A(_00931_),
    .B(_00986_),
    .C(_00953_),
    .Y(_01063_));
 sky130_fd_sc_hd__nand3_1 _15438_ (.A(_01019_),
    .B(_07713_),
    .C(_01008_),
    .Y(_01074_));
 sky130_fd_sc_hd__a21oi_4 _15439_ (.A1(_00855_),
    .A2(_00877_),
    .B1(_07713_),
    .Y(_01085_));
 sky130_fd_sc_hd__or3_1 _15440_ (.A(net372),
    .B(net371),
    .C(_00899_),
    .X(_01096_));
 sky130_fd_sc_hd__o221a_1 _15441_ (.A1(net372),
    .A2(net371),
    .B1(_00920_),
    .B2(_01052_),
    .C1(_01030_),
    .X(_01107_));
 sky130_fd_sc_hd__o221ai_4 _15442_ (.A1(net372),
    .A2(net371),
    .B1(_00920_),
    .B2(_01052_),
    .C1(_01030_),
    .Y(_01118_));
 sky130_fd_sc_hd__a31o_1 _15443_ (.A1(_01030_),
    .A2(_01063_),
    .A3(_07713_),
    .B1(_01085_),
    .X(_01129_));
 sky130_fd_sc_hd__a31o_1 _15444_ (.A1(_01019_),
    .A2(_07713_),
    .A3(_01008_),
    .B1(_00910_),
    .X(_01140_));
 sky130_fd_sc_hd__or4_1 _15445_ (.A(net353),
    .B(net352),
    .C(_01085_),
    .D(_01107_),
    .X(_01151_));
 sky130_fd_sc_hd__o32a_1 _15446_ (.A1(net380),
    .A2(net391),
    .A3(_13788_),
    .B1(_13832_),
    .B2(_13865_),
    .X(_01162_));
 sky130_fd_sc_hd__a311oi_4 _15447_ (.A1(_01030_),
    .A2(_01063_),
    .A3(_07713_),
    .B1(_01085_),
    .C1(_07044_),
    .Y(_01173_));
 sky130_fd_sc_hd__o221ai_4 _15448_ (.A1(_06989_),
    .A2(_07011_),
    .B1(_07713_),
    .B2(_00899_),
    .C1(_01118_),
    .Y(_01184_));
 sky130_fd_sc_hd__a2bb2oi_1 _15449_ (.A1_N(_06945_),
    .A2_N(net377),
    .B1(_01096_),
    .B2(_01118_),
    .Y(_01195_));
 sky130_fd_sc_hd__o211ai_4 _15450_ (.A1(_07713_),
    .A2(_00888_),
    .B1(_01074_),
    .C1(_07044_),
    .Y(_01206_));
 sky130_fd_sc_hd__o22ai_1 _15451_ (.A1(_13810_),
    .A2(_13909_),
    .B1(_01173_),
    .B2(_01195_),
    .Y(_01217_));
 sky130_fd_sc_hd__o2111ai_1 _15452_ (.A1(_06332_),
    .A2(_13788_),
    .B1(_13920_),
    .C1(_01184_),
    .D1(_01206_),
    .Y(_01228_));
 sky130_fd_sc_hd__nand3_2 _15453_ (.A(_01217_),
    .B(_01228_),
    .C(_08721_),
    .Y(_01239_));
 sky130_fd_sc_hd__a311o_1 _15454_ (.A1(_01019_),
    .A2(_07713_),
    .A3(_01008_),
    .B1(_08721_),
    .C1(_00910_),
    .X(_01250_));
 sky130_fd_sc_hd__o211ai_1 _15455_ (.A1(_13810_),
    .A2(_13909_),
    .B1(_01184_),
    .C1(_01206_),
    .Y(_01261_));
 sky130_fd_sc_hd__o21ai_1 _15456_ (.A1(_01173_),
    .A2(_01195_),
    .B1(_01162_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand3_1 _15457_ (.A(_01271_),
    .B(_08721_),
    .C(_01261_),
    .Y(_01282_));
 sky130_fd_sc_hd__o21ai_4 _15458_ (.A1(_08721_),
    .A2(_01129_),
    .B1(_01239_),
    .Y(_01293_));
 sky130_fd_sc_hd__o311a_4 _15459_ (.A1(_08721_),
    .A2(_01085_),
    .A3(_01107_),
    .B1(_01239_),
    .C1(_09840_),
    .X(_01304_));
 sky130_fd_sc_hd__inv_2 _15460_ (.A(_01304_),
    .Y(_01315_));
 sky130_fd_sc_hd__o211ai_2 _15461_ (.A1(net392),
    .A2(net382),
    .B1(_01151_),
    .C1(_01239_),
    .Y(_01326_));
 sky130_fd_sc_hd__o221a_1 _15462_ (.A1(net380),
    .A2(net391),
    .B1(_08721_),
    .B2(_01140_),
    .C1(_01282_),
    .X(_01337_));
 sky130_fd_sc_hd__nand3_1 _15463_ (.A(_01282_),
    .B(_06332_),
    .C(_01250_),
    .Y(_01348_));
 sky130_fd_sc_hd__a22oi_1 _15464_ (.A1(_13953_),
    .A2(_13975_),
    .B1(_14030_),
    .B2(_05862_),
    .Y(_01359_));
 sky130_fd_sc_hd__a21oi_1 _15465_ (.A1(_14129_),
    .A2(_14019_),
    .B1(_14140_),
    .Y(_01370_));
 sky130_fd_sc_hd__o32ai_4 _15466_ (.A1(_05862_),
    .A2(_13799_),
    .A3(_13931_),
    .B1(_14030_),
    .B2(_14118_),
    .Y(_01381_));
 sky130_fd_sc_hd__o2bb2ai_1 _15467_ (.A1_N(_01326_),
    .A2_N(_01348_),
    .B1(_01359_),
    .B2(_14041_),
    .Y(_01392_));
 sky130_fd_sc_hd__o211ai_2 _15468_ (.A1(_14030_),
    .A2(_14118_),
    .B1(_14151_),
    .C1(_01348_),
    .Y(_01403_));
 sky130_fd_sc_hd__nand3_1 _15469_ (.A(_01370_),
    .B(_01348_),
    .C(_01326_),
    .Y(_01414_));
 sky130_fd_sc_hd__and3_4 _15470_ (.A(_01392_),
    .B(_01414_),
    .C(_09829_),
    .X(_01425_));
 sky130_fd_sc_hd__nand3_2 _15471_ (.A(_01392_),
    .B(_01414_),
    .C(_09829_),
    .Y(_01436_));
 sky130_fd_sc_hd__a31o_1 _15472_ (.A1(_01392_),
    .A2(_01414_),
    .A3(_09829_),
    .B1(_01304_),
    .X(_01447_));
 sky130_fd_sc_hd__a31oi_2 _15473_ (.A1(_14184_),
    .A2(net385),
    .A3(_14107_),
    .B1(_14216_),
    .Y(_01458_));
 sky130_fd_sc_hd__o32ai_4 _15474_ (.A1(_05501_),
    .A2(_05523_),
    .A3(_14216_),
    .B1(_14227_),
    .B2(_14206_),
    .Y(_01469_));
 sky130_fd_sc_hd__o211ai_2 _15475_ (.A1(_14227_),
    .A2(_14206_),
    .B1(_05851_),
    .C1(_14249_),
    .Y(_01480_));
 sky130_fd_sc_hd__o22ai_4 _15476_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_14315_),
    .B2(_01458_),
    .Y(_01491_));
 sky130_fd_sc_hd__o311a_1 _15477_ (.A1(_05862_),
    .A2(_14315_),
    .A3(_01458_),
    .B1(_11068_),
    .C1(_01491_),
    .X(_01502_));
 sky130_fd_sc_hd__o2111ai_4 _15478_ (.A1(_01304_),
    .A2(_01425_),
    .B1(_11068_),
    .C1(_01480_),
    .D1(_01491_),
    .Y(_01513_));
 sky130_fd_sc_hd__a31o_1 _15479_ (.A1(_01491_),
    .A2(_11068_),
    .A3(_01480_),
    .B1(_01447_),
    .X(_01524_));
 sky130_fd_sc_hd__a211o_2 _15480_ (.A1(_01315_),
    .A2(_01436_),
    .B1(net347),
    .C1(net346),
    .X(_01535_));
 sky130_fd_sc_hd__a2bb2oi_4 _15481_ (.A1_N(_05763_),
    .A2_N(_05785_),
    .B1(_01315_),
    .B2(_01436_),
    .Y(_01546_));
 sky130_fd_sc_hd__o221a_1 _15482_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_09829_),
    .B2(_01293_),
    .C1(_01436_),
    .X(_01557_));
 sky130_fd_sc_hd__o21ai_1 _15483_ (.A1(_05862_),
    .A2(_01447_),
    .B1(_01469_),
    .Y(_01568_));
 sky130_fd_sc_hd__o21bai_1 _15484_ (.A1(_01546_),
    .A2(_01557_),
    .B1_N(_01469_),
    .Y(_01579_));
 sky130_fd_sc_hd__o221ai_4 _15485_ (.A1(net347),
    .A2(net346),
    .B1(_01546_),
    .B2(_01568_),
    .C1(_01579_),
    .Y(_01590_));
 sky130_fd_sc_hd__nand2_2 _15486_ (.A(_01535_),
    .B(_01590_),
    .Y(_01600_));
 sky130_fd_sc_hd__o32a_1 _15487_ (.A1(_05250_),
    .A2(_14271_),
    .A3(_14293_),
    .B1(_12637_),
    .B2(_14348_),
    .X(_01611_));
 sky130_fd_sc_hd__o32ai_4 _15488_ (.A1(_05250_),
    .A2(_14271_),
    .A3(_14293_),
    .B1(_12637_),
    .B2(_14348_),
    .Y(_01622_));
 sky130_fd_sc_hd__o221ai_4 _15489_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_12637_),
    .B2(_14348_),
    .C1(_14337_),
    .Y(_01633_));
 sky130_fd_sc_hd__o21ai_4 _15490_ (.A1(net398),
    .A2(net397),
    .B1(_01622_),
    .Y(_01644_));
 sky130_fd_sc_hd__o2111a_1 _15491_ (.A1(net328),
    .A2(_12681_),
    .B1(_01600_),
    .C1(_01633_),
    .D1(_01644_),
    .X(_01655_));
 sky130_fd_sc_hd__o2111ai_4 _15492_ (.A1(net328),
    .A2(_12681_),
    .B1(_01600_),
    .C1(_01633_),
    .D1(_01644_),
    .Y(_01666_));
 sky130_fd_sc_hd__a31oi_4 _15493_ (.A1(_01644_),
    .A2(_12692_),
    .A3(_01633_),
    .B1(_01600_),
    .Y(_01677_));
 sky130_fd_sc_hd__a31o_1 _15494_ (.A1(_01644_),
    .A2(_12692_),
    .A3(_01633_),
    .B1(_01600_),
    .X(_01688_));
 sky130_fd_sc_hd__nand3_1 _15495_ (.A(_01590_),
    .B(net385),
    .C(_01535_),
    .Y(_01699_));
 sky130_fd_sc_hd__o211a_2 _15496_ (.A1(net398),
    .A2(net397),
    .B1(_01513_),
    .C1(_01524_),
    .X(_01710_));
 sky130_fd_sc_hd__o211ai_4 _15497_ (.A1(net398),
    .A2(net397),
    .B1(_01513_),
    .C1(_01524_),
    .Y(_01721_));
 sky130_fd_sc_hd__nand3_1 _15498_ (.A(_01622_),
    .B(_01699_),
    .C(_01721_),
    .Y(_01732_));
 sky130_fd_sc_hd__a21o_1 _15499_ (.A1(_01699_),
    .A2(_01721_),
    .B1(_01622_),
    .X(_01743_));
 sky130_fd_sc_hd__nand3_1 _15500_ (.A(_01743_),
    .B(_12692_),
    .C(_01732_),
    .Y(_01754_));
 sky130_fd_sc_hd__o311a_1 _15501_ (.A1(_01304_),
    .A2(_01425_),
    .A3(_01502_),
    .B1(_01513_),
    .C1(_12703_),
    .X(_01765_));
 sky130_fd_sc_hd__a211o_1 _15502_ (.A1(_01535_),
    .A2(_01590_),
    .B1(net328),
    .C1(_12681_),
    .X(_01776_));
 sky130_fd_sc_hd__nor3_2 _15503_ (.A(_05250_),
    .B(_01655_),
    .C(_01677_),
    .Y(_01787_));
 sky130_fd_sc_hd__nand3_4 _15504_ (.A(_01688_),
    .B(net403),
    .C(_01666_),
    .Y(_01798_));
 sky130_fd_sc_hd__a311oi_4 _15505_ (.A1(_01743_),
    .A2(_12692_),
    .A3(_01732_),
    .B1(_01765_),
    .C1(net403),
    .Y(_01809_));
 sky130_fd_sc_hd__o21ai_2 _15506_ (.A1(_01655_),
    .A2(_01677_),
    .B1(_05250_),
    .Y(_01820_));
 sky130_fd_sc_hd__o41a_1 _15507_ (.A1(_05196_),
    .A2(_05218_),
    .A3(_01655_),
    .A4(_01677_),
    .B1(_01820_),
    .X(_01831_));
 sky130_fd_sc_hd__a31oi_2 _15508_ (.A1(_05250_),
    .A2(_01754_),
    .A3(_01776_),
    .B1(_14425_),
    .Y(_01842_));
 sky130_fd_sc_hd__nand2_1 _15509_ (.A(_01820_),
    .B(_14414_),
    .Y(_01853_));
 sky130_fd_sc_hd__a31oi_1 _15510_ (.A1(_01820_),
    .A2(_14414_),
    .A3(_01798_),
    .B1(_00066_),
    .Y(_01864_));
 sky130_fd_sc_hd__o21ai_1 _15511_ (.A1(_14414_),
    .A2(_01831_),
    .B1(_01864_),
    .Y(_01875_));
 sky130_fd_sc_hd__or4_1 _15512_ (.A(net324),
    .B(net322),
    .C(_01655_),
    .D(_01677_),
    .X(_01886_));
 sky130_fd_sc_hd__nand2_1 _15513_ (.A(_01875_),
    .B(_01886_),
    .Y(_01897_));
 sky130_fd_sc_hd__or3_4 _15514_ (.A(net64),
    .B(net34),
    .C(_12659_),
    .X(_01908_));
 sky130_fd_sc_hd__o311a_4 _15515_ (.A1(net64),
    .A2(net34),
    .A3(_12659_),
    .B1(net35),
    .C1(net409),
    .X(_01919_));
 sky130_fd_sc_hd__a21oi_4 _15516_ (.A1(_01908_),
    .A2(net409),
    .B1(net35),
    .Y(_01930_));
 sky130_fd_sc_hd__a21boi_4 _15517_ (.A1(_01908_),
    .A2(net409),
    .B1_N(net35),
    .Y(_01940_));
 sky130_fd_sc_hd__and3b_4 _15518_ (.A_N(net35),
    .B(_01908_),
    .C(net409),
    .X(_01951_));
 sky130_fd_sc_hd__nor2_8 _15519_ (.A(_01919_),
    .B(_01930_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_8 _15520_ (.A(net304),
    .B(_01951_),
    .Y(_01973_));
 sky130_fd_sc_hd__o311a_1 _15521_ (.A1(_03289_),
    .A2(_01919_),
    .A3(_01930_),
    .B1(_01875_),
    .C1(_01886_),
    .X(_01984_));
 sky130_fd_sc_hd__a21oi_1 _15522_ (.A1(_01875_),
    .A2(_01886_),
    .B1(_03289_),
    .Y(_01995_));
 sky130_fd_sc_hd__a31oi_1 _15523_ (.A1(net1),
    .A2(_01897_),
    .A3(_01962_),
    .B1(_01984_),
    .Y(_02006_));
 sky130_fd_sc_hd__xnor2_1 _15524_ (.A(_00109_),
    .B(_02006_),
    .Y(net67));
 sky130_fd_sc_hd__and3b_1 _15525_ (.A_N(_02006_),
    .B(_00088_),
    .C(_12746_),
    .X(_02027_));
 sky130_fd_sc_hd__or4_4 _15526_ (.A(net2),
    .B(_12823_),
    .C(net3),
    .D(_09916_),
    .X(_02038_));
 sky130_fd_sc_hd__and3_4 _15527_ (.A(_02038_),
    .B(net410),
    .C(_04503_),
    .X(_02049_));
 sky130_fd_sc_hd__a311o_4 _15528_ (.A1(_12834_),
    .A2(_04392_),
    .A3(_04282_),
    .B1(_03399_),
    .C1(net4),
    .X(_02060_));
 sky130_fd_sc_hd__a21oi_4 _15529_ (.A1(_02038_),
    .A2(net410),
    .B1(_04503_),
    .Y(_02071_));
 sky130_fd_sc_hd__a21o_4 _15530_ (.A1(_02038_),
    .A2(net410),
    .B1(_04503_),
    .X(_02082_));
 sky130_fd_sc_hd__a21oi_4 _15531_ (.A1(_02038_),
    .A2(net410),
    .B1(net4),
    .Y(_02093_));
 sky130_fd_sc_hd__a21o_4 _15532_ (.A1(_02038_),
    .A2(net410),
    .B1(net4),
    .X(_02104_));
 sky130_fd_sc_hd__and3_4 _15533_ (.A(_02038_),
    .B(net4),
    .C(net410),
    .X(_02115_));
 sky130_fd_sc_hd__a311o_4 _15534_ (.A1(_12834_),
    .A2(_04392_),
    .A3(_04282_),
    .B1(_03399_),
    .C1(_04503_),
    .X(_02126_));
 sky130_fd_sc_hd__nand2_8 _15535_ (.A(_02104_),
    .B(_02126_),
    .Y(_02137_));
 sky130_fd_sc_hd__nand2_8 _15536_ (.A(_02060_),
    .B(_02082_),
    .Y(_02148_));
 sky130_fd_sc_hd__or3_2 _15537_ (.A(_03178_),
    .B(_02093_),
    .C(_02115_),
    .X(_02159_));
 sky130_fd_sc_hd__o221a_1 _15538_ (.A1(net408),
    .A2(_05152_),
    .B1(_02049_),
    .B2(net342),
    .C1(net33),
    .X(_02170_));
 sky130_fd_sc_hd__or4_1 _15539_ (.A(_03178_),
    .B(_05174_),
    .C(_02093_),
    .D(_02115_),
    .X(_02181_));
 sky130_fd_sc_hd__a31o_1 _15540_ (.A1(_02104_),
    .A2(_02126_),
    .A3(net33),
    .B1(net319),
    .X(_02192_));
 sky130_fd_sc_hd__o31a_1 _15541_ (.A1(_00273_),
    .A2(_02093_),
    .A3(_02115_),
    .B1(_02192_),
    .X(_02203_));
 sky130_fd_sc_hd__o21ai_2 _15542_ (.A1(_00273_),
    .A2(_02137_),
    .B1(_02192_),
    .Y(_02214_));
 sky130_fd_sc_hd__o211ai_2 _15543_ (.A1(net320),
    .A2(_12910_),
    .B1(_12932_),
    .C1(_13075_),
    .Y(_02225_));
 sky130_fd_sc_hd__o221ai_4 _15544_ (.A1(_12910_),
    .A2(net320),
    .B1(_00306_),
    .B2(_00284_),
    .C1(_02214_),
    .Y(_02236_));
 sky130_fd_sc_hd__o211ai_4 _15545_ (.A1(net325),
    .A2(_00262_),
    .B1(_02203_),
    .C1(_02225_),
    .Y(_02247_));
 sky130_fd_sc_hd__nand2_1 _15546_ (.A(_02236_),
    .B(_02247_),
    .Y(_02258_));
 sky130_fd_sc_hd__nand3_1 _15547_ (.A(_02236_),
    .B(_02247_),
    .C(_05174_),
    .Y(_02268_));
 sky130_fd_sc_hd__o32a_1 _15548_ (.A1(_03178_),
    .A2(_02093_),
    .A3(_02115_),
    .B1(net408),
    .B2(_05152_),
    .X(_02279_));
 sky130_fd_sc_hd__a31o_1 _15549_ (.A1(_02104_),
    .A2(_02126_),
    .A3(net33),
    .B1(_05174_),
    .X(_02290_));
 sky130_fd_sc_hd__o31a_1 _15550_ (.A1(_03178_),
    .A2(_05174_),
    .A3(_02137_),
    .B1(_02268_),
    .X(_02301_));
 sky130_fd_sc_hd__a31o_1 _15551_ (.A1(_02236_),
    .A2(_02247_),
    .A3(_05174_),
    .B1(_02170_),
    .X(_02312_));
 sky130_fd_sc_hd__and3_1 _15552_ (.A(_05359_),
    .B(_05381_),
    .C(_02312_),
    .X(_02323_));
 sky130_fd_sc_hd__or3_4 _15553_ (.A(net402),
    .B(net400),
    .C(_02301_),
    .X(_02334_));
 sky130_fd_sc_hd__o311a_2 _15554_ (.A1(_03178_),
    .A2(_05174_),
    .A3(_02137_),
    .B1(_12888_),
    .C1(_02268_),
    .X(_02345_));
 sky130_fd_sc_hd__a311o_4 _15555_ (.A1(_02236_),
    .A2(_02247_),
    .A3(_05174_),
    .B1(net325),
    .C1(_02170_),
    .X(_02356_));
 sky130_fd_sc_hd__o2bb2a_1 _15556_ (.A1_N(_05174_),
    .A2_N(_02258_),
    .B1(_12856_),
    .B2(_12845_),
    .X(_02367_));
 sky130_fd_sc_hd__a2bb2o_1 _15557_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_05174_),
    .B2(_02258_),
    .X(_02378_));
 sky130_fd_sc_hd__a21oi_1 _15558_ (.A1(_02181_),
    .A2(_02268_),
    .B1(_12888_),
    .Y(_02389_));
 sky130_fd_sc_hd__o21ai_2 _15559_ (.A1(_12845_),
    .A2(_12856_),
    .B1(_02312_),
    .Y(_02400_));
 sky130_fd_sc_hd__nor2_1 _15560_ (.A(_02345_),
    .B(_02389_),
    .Y(_02411_));
 sky130_fd_sc_hd__nand2_1 _15561_ (.A(_02356_),
    .B(_02400_),
    .Y(_02422_));
 sky130_fd_sc_hd__a31oi_4 _15562_ (.A1(_13185_),
    .A2(_00438_),
    .A3(_00482_),
    .B1(_00449_),
    .Y(_02433_));
 sky130_fd_sc_hd__a31o_1 _15563_ (.A1(_13185_),
    .A2(_00438_),
    .A3(_00482_),
    .B1(_00449_),
    .X(_02444_));
 sky130_fd_sc_hd__o21ai_2 _15564_ (.A1(_02345_),
    .A2(_02389_),
    .B1(_02433_),
    .Y(_02455_));
 sky130_fd_sc_hd__a22oi_2 _15565_ (.A1(_05359_),
    .A2(_05381_),
    .B1(_02411_),
    .B2(_02444_),
    .Y(_02466_));
 sky130_fd_sc_hd__o211a_1 _15566_ (.A1(_02433_),
    .A2(_02422_),
    .B1(net388),
    .C1(_02455_),
    .X(_02477_));
 sky130_fd_sc_hd__o211ai_4 _15567_ (.A1(_02433_),
    .A2(_02422_),
    .B1(net388),
    .C1(_02455_),
    .Y(_02488_));
 sky130_fd_sc_hd__a22o_2 _15568_ (.A1(_05392_),
    .A2(_02312_),
    .B1(_02466_),
    .B2(_02455_),
    .X(_02499_));
 sky130_fd_sc_hd__and3_1 _15569_ (.A(_05687_),
    .B(_05709_),
    .C(_02499_),
    .X(_02510_));
 sky130_fd_sc_hd__a211o_2 _15570_ (.A1(_02334_),
    .A2(_02488_),
    .B1(net384),
    .C1(net383),
    .X(_02521_));
 sky130_fd_sc_hd__a2bb2oi_4 _15571_ (.A1_N(_11210_),
    .A2_N(_11232_),
    .B1(_02334_),
    .B2(_02488_),
    .Y(_02532_));
 sky130_fd_sc_hd__o22ai_4 _15572_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_02323_),
    .B2(_02477_),
    .Y(_02543_));
 sky130_fd_sc_hd__a22oi_2 _15573_ (.A1(_11265_),
    .A2(_11287_),
    .B1(_02466_),
    .B2(_02455_),
    .Y(_02554_));
 sky130_fd_sc_hd__o21ai_1 _15574_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_02488_),
    .Y(_02564_));
 sky130_fd_sc_hd__o211a_1 _15575_ (.A1(net388),
    .A2(_02301_),
    .B1(net331),
    .C1(_02488_),
    .X(_02575_));
 sky130_fd_sc_hd__o211ai_4 _15576_ (.A1(net388),
    .A2(_02301_),
    .B1(net331),
    .C1(_02488_),
    .Y(_02586_));
 sky130_fd_sc_hd__a31oi_2 _15577_ (.A1(_13415_),
    .A2(_00646_),
    .A3(_00657_),
    .B1(_00613_),
    .Y(_02597_));
 sky130_fd_sc_hd__o41ai_4 _15578_ (.A1(_09971_),
    .A2(net363),
    .A3(_00547_),
    .A4(_00558_),
    .B1(_00745_),
    .Y(_02608_));
 sky130_fd_sc_hd__a221oi_4 _15579_ (.A1(_02554_),
    .A2(_02334_),
    .B1(_00745_),
    .B2(_00624_),
    .C1(_02532_),
    .Y(_02619_));
 sky130_fd_sc_hd__o211ai_2 _15580_ (.A1(_02564_),
    .A2(_02323_),
    .B1(_02543_),
    .C1(_02608_),
    .Y(_02630_));
 sky130_fd_sc_hd__a21oi_2 _15581_ (.A1(_02543_),
    .A2(_02586_),
    .B1(_02608_),
    .Y(_02641_));
 sky130_fd_sc_hd__o21ai_2 _15582_ (.A1(_02532_),
    .A2(_02575_),
    .B1(_02597_),
    .Y(_02652_));
 sky130_fd_sc_hd__nand3_4 _15583_ (.A(_02652_),
    .B(_05720_),
    .C(_02630_),
    .Y(_02663_));
 sky130_fd_sc_hd__o22ai_4 _15584_ (.A1(net384),
    .A2(net383),
    .B1(_02619_),
    .B2(_02641_),
    .Y(_02674_));
 sky130_fd_sc_hd__a2bb2oi_4 _15585_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_02521_),
    .B2(_02663_),
    .Y(_02685_));
 sky130_fd_sc_hd__o211ai_4 _15586_ (.A1(_02499_),
    .A2(_05720_),
    .B1(net348),
    .C1(_02674_),
    .Y(_02696_));
 sky130_fd_sc_hd__o32a_4 _15587_ (.A1(_08863_),
    .A2(net366),
    .A3(_00778_),
    .B1(_00789_),
    .B2(_00142_),
    .X(_02707_));
 sky130_fd_sc_hd__o32ai_4 _15588_ (.A1(_08863_),
    .A2(net366),
    .A3(_00778_),
    .B1(_00789_),
    .B2(_00142_),
    .Y(_02718_));
 sky130_fd_sc_hd__a31o_1 _15589_ (.A1(_02652_),
    .A2(_05720_),
    .A3(_02630_),
    .B1(net348),
    .X(_02729_));
 sky130_fd_sc_hd__o211a_1 _15590_ (.A1(_09971_),
    .A2(net363),
    .B1(_02521_),
    .C1(_02663_),
    .X(_02740_));
 sky130_fd_sc_hd__o211ai_4 _15591_ (.A1(_09971_),
    .A2(net363),
    .B1(_02521_),
    .C1(_02663_),
    .Y(_02751_));
 sky130_fd_sc_hd__o21ai_1 _15592_ (.A1(_02510_),
    .A2(_02729_),
    .B1(_02718_),
    .Y(_02762_));
 sky130_fd_sc_hd__nand3_4 _15593_ (.A(_02696_),
    .B(_02718_),
    .C(_02751_),
    .Y(_02773_));
 sky130_fd_sc_hd__o21ai_4 _15594_ (.A1(_02685_),
    .A2(_02740_),
    .B1(_02707_),
    .Y(_02784_));
 sky130_fd_sc_hd__and3_1 _15595_ (.A(_02784_),
    .B(_06837_),
    .C(_02773_),
    .X(_02795_));
 sky130_fd_sc_hd__nand3_2 _15596_ (.A(_02784_),
    .B(_06837_),
    .C(_02773_),
    .Y(_02806_));
 sky130_fd_sc_hd__o311a_4 _15597_ (.A1(net384),
    .A2(_02499_),
    .A3(net383),
    .B1(_06848_),
    .C1(_02674_),
    .X(_02817_));
 sky130_fd_sc_hd__a211o_1 _15598_ (.A1(_02521_),
    .A2(_02663_),
    .B1(net379),
    .C1(net378),
    .X(_02828_));
 sky130_fd_sc_hd__o311a_2 _15599_ (.A1(_05731_),
    .A2(_02619_),
    .A3(_02641_),
    .B1(_06848_),
    .C1(_02521_),
    .X(_02839_));
 sky130_fd_sc_hd__a21oi_1 _15600_ (.A1(_02773_),
    .A2(_02784_),
    .B1(_06848_),
    .Y(_02850_));
 sky130_fd_sc_hd__a31oi_4 _15601_ (.A1(_13679_),
    .A2(_00953_),
    .A3(_00964_),
    .B1(_00920_),
    .Y(_02860_));
 sky130_fd_sc_hd__o21ai_1 _15602_ (.A1(_07888_),
    .A2(_00899_),
    .B1(_01052_),
    .Y(_02871_));
 sky130_fd_sc_hd__o22ai_2 _15603_ (.A1(_08819_),
    .A2(net367),
    .B1(_00920_),
    .B2(_01041_),
    .Y(_02882_));
 sky130_fd_sc_hd__a31oi_4 _15604_ (.A1(_01052_),
    .A2(_08907_),
    .A3(_00931_),
    .B1(_07724_),
    .Y(_02893_));
 sky130_fd_sc_hd__o2bb2ai_4 _15605_ (.A1_N(_02882_),
    .A2_N(_02893_),
    .B1(_02839_),
    .B2(_02850_),
    .Y(_02904_));
 sky130_fd_sc_hd__o221ai_4 _15606_ (.A1(_02795_),
    .A2(_02817_),
    .B1(_02860_),
    .B2(_08907_),
    .C1(_02893_),
    .Y(_02915_));
 sky130_fd_sc_hd__or4_1 _15607_ (.A(net372),
    .B(net371),
    .C(_02839_),
    .D(_02850_),
    .X(_02926_));
 sky130_fd_sc_hd__a31o_1 _15608_ (.A1(_02784_),
    .A2(_06837_),
    .A3(_02773_),
    .B1(_08918_),
    .X(_02937_));
 sky130_fd_sc_hd__a311oi_4 _15609_ (.A1(_02784_),
    .A2(_06837_),
    .A3(_02773_),
    .B1(_02817_),
    .C1(_08918_),
    .Y(_02948_));
 sky130_fd_sc_hd__a22oi_4 _15610_ (.A1(_08830_),
    .A2(_08852_),
    .B1(_02806_),
    .B2(_02828_),
    .Y(_02959_));
 sky130_fd_sc_hd__a22o_1 _15611_ (.A1(_08830_),
    .A2(_08852_),
    .B1(_02806_),
    .B2(_02828_),
    .X(_02970_));
 sky130_fd_sc_hd__o221ai_1 _15612_ (.A1(_00920_),
    .A2(_01041_),
    .B1(_02817_),
    .B2(_02937_),
    .C1(_02970_),
    .Y(_02981_));
 sky130_fd_sc_hd__o21ai_1 _15613_ (.A1(_02948_),
    .A2(_02959_),
    .B1(_02860_),
    .Y(_02992_));
 sky130_fd_sc_hd__nand3_1 _15614_ (.A(_02992_),
    .B(_07713_),
    .C(_02981_),
    .Y(_03003_));
 sky130_fd_sc_hd__nand2_1 _15615_ (.A(_02926_),
    .B(_03003_),
    .Y(_03014_));
 sky130_fd_sc_hd__o311a_1 _15616_ (.A1(net380),
    .A2(net391),
    .A3(_13788_),
    .B1(_13920_),
    .C1(_01206_),
    .X(_03025_));
 sky130_fd_sc_hd__o211ai_2 _15617_ (.A1(_06332_),
    .A2(_13788_),
    .B1(_13920_),
    .C1(_01206_),
    .Y(_03036_));
 sky130_fd_sc_hd__o2bb2ai_2 _15618_ (.A1_N(_13821_),
    .A2_N(_13920_),
    .B1(_07044_),
    .B2(_01129_),
    .Y(_03047_));
 sky130_fd_sc_hd__a21oi_4 _15619_ (.A1(_02904_),
    .A2(_02915_),
    .B1(_07899_),
    .Y(_03058_));
 sky130_fd_sc_hd__nand3_2 _15620_ (.A(_03003_),
    .B(_07888_),
    .C(_02926_),
    .Y(_03069_));
 sky130_fd_sc_hd__o211a_1 _15621_ (.A1(net389),
    .A2(net370),
    .B1(_02904_),
    .C1(_02915_),
    .X(_03080_));
 sky130_fd_sc_hd__nand3_4 _15622_ (.A(_07899_),
    .B(_02904_),
    .C(_02915_),
    .Y(_03091_));
 sky130_fd_sc_hd__o311a_1 _15623_ (.A1(_07044_),
    .A2(_01085_),
    .A3(_01107_),
    .B1(_03036_),
    .C1(_03069_),
    .X(_03102_));
 sky130_fd_sc_hd__nand4_4 _15624_ (.A(_01184_),
    .B(_03036_),
    .C(_03069_),
    .D(_03091_),
    .Y(_03113_));
 sky130_fd_sc_hd__o22ai_4 _15625_ (.A1(_01173_),
    .A2(_03025_),
    .B1(_03058_),
    .B2(_03080_),
    .Y(_03123_));
 sky130_fd_sc_hd__and3_2 _15626_ (.A(_08732_),
    .B(_02904_),
    .C(_02915_),
    .X(_03134_));
 sky130_fd_sc_hd__a211o_2 _15627_ (.A1(_02926_),
    .A2(_03003_),
    .B1(net353),
    .C1(net352),
    .X(_03145_));
 sky130_fd_sc_hd__nand3_2 _15628_ (.A(_03123_),
    .B(_08721_),
    .C(_03113_),
    .Y(_03156_));
 sky130_fd_sc_hd__a31o_1 _15629_ (.A1(_03123_),
    .A2(_08721_),
    .A3(_03113_),
    .B1(_03134_),
    .X(_03167_));
 sky130_fd_sc_hd__a31oi_4 _15630_ (.A1(_03123_),
    .A2(_08721_),
    .A3(_03113_),
    .B1(_03134_),
    .Y(_03179_));
 sky130_fd_sc_hd__and3_1 _15631_ (.A(_03167_),
    .B(_09818_),
    .C(_09796_),
    .X(_03190_));
 sky130_fd_sc_hd__or3_1 _15632_ (.A(net350),
    .B(net349),
    .C(_03179_),
    .X(_03201_));
 sky130_fd_sc_hd__o32a_1 _15633_ (.A1(net380),
    .A2(net391),
    .A3(_01293_),
    .B1(_01381_),
    .B2(_01337_),
    .X(_03212_));
 sky130_fd_sc_hd__o32ai_4 _15634_ (.A1(net380),
    .A2(net391),
    .A3(_01293_),
    .B1(_01381_),
    .B2(_01337_),
    .Y(_03223_));
 sky130_fd_sc_hd__a311oi_4 _15635_ (.A1(_03123_),
    .A2(_08721_),
    .A3(_03113_),
    .B1(_03134_),
    .C1(_07044_),
    .Y(_03234_));
 sky130_fd_sc_hd__o211ai_4 _15636_ (.A1(_06989_),
    .A2(_07011_),
    .B1(_03145_),
    .C1(_03156_),
    .Y(_03245_));
 sky130_fd_sc_hd__a2bb2oi_2 _15637_ (.A1_N(_06945_),
    .A2_N(net377),
    .B1(_03145_),
    .B2(_03156_),
    .Y(_03256_));
 sky130_fd_sc_hd__a22o_1 _15638_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_03145_),
    .B2(_03156_),
    .X(_03267_));
 sky130_fd_sc_hd__o2bb2ai_1 _15639_ (.A1_N(_01326_),
    .A2_N(_01403_),
    .B1(_03179_),
    .B2(_07033_),
    .Y(_03278_));
 sky130_fd_sc_hd__nand3_2 _15640_ (.A(_03223_),
    .B(_03245_),
    .C(_03267_),
    .Y(_03290_));
 sky130_fd_sc_hd__o21ai_4 _15641_ (.A1(_03234_),
    .A2(_03256_),
    .B1(_03212_),
    .Y(_03301_));
 sky130_fd_sc_hd__o211ai_4 _15642_ (.A1(_03234_),
    .A2(_03278_),
    .B1(_09829_),
    .C1(_03301_),
    .Y(_03312_));
 sky130_fd_sc_hd__a31oi_4 _15643_ (.A1(_03290_),
    .A2(_03301_),
    .A3(net337),
    .B1(_03190_),
    .Y(_03323_));
 sky130_fd_sc_hd__inv_2 _15644_ (.A(_03323_),
    .Y(_03334_));
 sky130_fd_sc_hd__or3_2 _15645_ (.A(net347),
    .B(net346),
    .C(_03323_),
    .X(_03345_));
 sky130_fd_sc_hd__a2bb2oi_1 _15646_ (.A1_N(net392),
    .A2_N(net382),
    .B1(_03201_),
    .B2(_03312_),
    .Y(_03356_));
 sky130_fd_sc_hd__a22o_1 _15647_ (.A1(_06256_),
    .A2(_06278_),
    .B1(_03201_),
    .B2(_03312_),
    .X(_03367_));
 sky130_fd_sc_hd__o221a_2 _15648_ (.A1(net380),
    .A2(net391),
    .B1(_09829_),
    .B2(_03179_),
    .C1(_03312_),
    .X(_03378_));
 sky130_fd_sc_hd__o221ai_4 _15649_ (.A1(net380),
    .A2(net391),
    .B1(_09829_),
    .B2(_03179_),
    .C1(_03312_),
    .Y(_03388_));
 sky130_fd_sc_hd__o32a_1 _15650_ (.A1(_05862_),
    .A2(_01304_),
    .A3(_01425_),
    .B1(_01469_),
    .B2(_01546_),
    .X(_03400_));
 sky130_fd_sc_hd__o32ai_4 _15651_ (.A1(_05862_),
    .A2(_01304_),
    .A3(_01425_),
    .B1(_01469_),
    .B2(_01546_),
    .Y(_03411_));
 sky130_fd_sc_hd__o21ai_1 _15652_ (.A1(_03356_),
    .A2(_03378_),
    .B1(_03400_),
    .Y(_03422_));
 sky130_fd_sc_hd__nand3_1 _15653_ (.A(_03367_),
    .B(_03388_),
    .C(_03411_),
    .Y(_03433_));
 sky130_fd_sc_hd__o21ai_1 _15654_ (.A1(_03356_),
    .A2(_03378_),
    .B1(_03411_),
    .Y(_03444_));
 sky130_fd_sc_hd__nand3_1 _15655_ (.A(_03367_),
    .B(_03388_),
    .C(_03400_),
    .Y(_03455_));
 sky130_fd_sc_hd__nand3_1 _15656_ (.A(_03444_),
    .B(_03455_),
    .C(_11068_),
    .Y(_03466_));
 sky130_fd_sc_hd__nand3_2 _15657_ (.A(_03422_),
    .B(_03433_),
    .C(_11068_),
    .Y(_03477_));
 sky130_fd_sc_hd__a311o_1 _15658_ (.A1(_03290_),
    .A2(_03301_),
    .A3(net337),
    .B1(_11068_),
    .C1(_03190_),
    .X(_03488_));
 sky130_fd_sc_hd__o31a_2 _15659_ (.A1(net347),
    .A2(net346),
    .A3(_03334_),
    .B1(_03477_),
    .X(_03499_));
 sky130_fd_sc_hd__o311ai_4 _15660_ (.A1(_01304_),
    .A2(_01425_),
    .A3(_01502_),
    .B1(_01513_),
    .C1(_01622_),
    .Y(_03511_));
 sky130_fd_sc_hd__a32oi_4 _15661_ (.A1(_01590_),
    .A2(net385),
    .A3(_01535_),
    .B1(_14337_),
    .B2(_14381_),
    .Y(_03522_));
 sky130_fd_sc_hd__a21oi_2 _15662_ (.A1(_01622_),
    .A2(_01699_),
    .B1(_01710_),
    .Y(_03533_));
 sky130_fd_sc_hd__a32o_1 _15663_ (.A1(_05512_),
    .A2(_05534_),
    .A3(_01622_),
    .B1(_01600_),
    .B2(_01633_),
    .X(_03544_));
 sky130_fd_sc_hd__o2111ai_4 _15664_ (.A1(net385),
    .A2(_01611_),
    .B1(_01721_),
    .C1(_05851_),
    .D1(_03511_),
    .Y(_03555_));
 sky130_fd_sc_hd__o22ai_4 _15665_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_01710_),
    .B2(_03522_),
    .Y(_03566_));
 sky130_fd_sc_hd__o311a_1 _15666_ (.A1(_05862_),
    .A2(_01710_),
    .A3(_03522_),
    .B1(_12692_),
    .C1(_03566_),
    .X(_03577_));
 sky130_fd_sc_hd__a31oi_2 _15667_ (.A1(_03566_),
    .A2(_12692_),
    .A3(_03555_),
    .B1(_03499_),
    .Y(_03588_));
 sky130_fd_sc_hd__a31o_1 _15668_ (.A1(_03566_),
    .A2(_12692_),
    .A3(_03555_),
    .B1(_03499_),
    .X(_03599_));
 sky130_fd_sc_hd__nand4_4 _15669_ (.A(_03499_),
    .B(_03555_),
    .C(_03566_),
    .D(_12692_),
    .Y(_03610_));
 sky130_fd_sc_hd__a211o_1 _15670_ (.A1(_03345_),
    .A2(_03466_),
    .B1(net328),
    .C1(_12681_),
    .X(_03622_));
 sky130_fd_sc_hd__o211ai_4 _15671_ (.A1(_03334_),
    .A2(_11068_),
    .B1(_05862_),
    .C1(_03477_),
    .Y(_03632_));
 sky130_fd_sc_hd__a31oi_2 _15672_ (.A1(_03444_),
    .A2(_03455_),
    .A3(_11068_),
    .B1(_05862_),
    .Y(_03643_));
 sky130_fd_sc_hd__nand3_1 _15673_ (.A(_03466_),
    .B(_05851_),
    .C(_03345_),
    .Y(_03654_));
 sky130_fd_sc_hd__o211ai_1 _15674_ (.A1(_03522_),
    .A2(_01710_),
    .B1(_03654_),
    .C1(_03632_),
    .Y(_03665_));
 sky130_fd_sc_hd__a21o_1 _15675_ (.A1(_03632_),
    .A2(_03654_),
    .B1(_03544_),
    .X(_03676_));
 sky130_fd_sc_hd__o211ai_1 _15676_ (.A1(net328),
    .A2(_12681_),
    .B1(_03665_),
    .C1(_03676_),
    .Y(_03687_));
 sky130_fd_sc_hd__a31oi_4 _15677_ (.A1(_03577_),
    .A2(_03488_),
    .A3(_03477_),
    .B1(_03588_),
    .Y(_03698_));
 sky130_fd_sc_hd__nand2_2 _15678_ (.A(_03599_),
    .B(_03610_),
    .Y(_03709_));
 sky130_fd_sc_hd__a21oi_4 _15679_ (.A1(_01820_),
    .A2(_14414_),
    .B1(_01787_),
    .Y(_03720_));
 sky130_fd_sc_hd__o21ai_2 _15680_ (.A1(_14425_),
    .A2(_01809_),
    .B1(_01798_),
    .Y(_03732_));
 sky130_fd_sc_hd__o221ai_4 _15681_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_14425_),
    .B2(_01809_),
    .C1(_01798_),
    .Y(_03743_));
 sky130_fd_sc_hd__a2bb2oi_2 _15682_ (.A1_N(net398),
    .A2_N(net397),
    .B1(_01798_),
    .B2(_01853_),
    .Y(_03754_));
 sky130_fd_sc_hd__o22ai_4 _15683_ (.A1(net398),
    .A2(net397),
    .B1(_01787_),
    .B2(_01842_),
    .Y(_03765_));
 sky130_fd_sc_hd__and4_1 _15684_ (.A(_03765_),
    .B(_00055_),
    .C(_03743_),
    .D(_03698_),
    .X(_03776_));
 sky130_fd_sc_hd__o2111ai_4 _15685_ (.A1(net324),
    .A2(net322),
    .B1(_03698_),
    .C1(_03743_),
    .D1(_03765_),
    .Y(_03787_));
 sky130_fd_sc_hd__a31oi_2 _15686_ (.A1(_03765_),
    .A2(_00055_),
    .A3(_03743_),
    .B1(_03698_),
    .Y(_03798_));
 sky130_fd_sc_hd__a31o_1 _15687_ (.A1(_03765_),
    .A2(_00055_),
    .A3(_03743_),
    .B1(_03698_),
    .X(_03809_));
 sky130_fd_sc_hd__o211ai_2 _15688_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_03622_),
    .C1(_03687_),
    .Y(_03820_));
 sky130_fd_sc_hd__o2111ai_4 _15689_ (.A1(_03399_),
    .A2(_05491_),
    .B1(_05534_),
    .C1(_03599_),
    .D1(_03610_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand4_1 _15690_ (.A(_05207_),
    .B(_05229_),
    .C(_03787_),
    .D(_03809_),
    .Y(_03842_));
 sky130_fd_sc_hd__a21oi_1 _15691_ (.A1(_03787_),
    .A2(_03809_),
    .B1(net403),
    .Y(_03853_));
 sky130_fd_sc_hd__o21ai_4 _15692_ (.A1(_03776_),
    .A2(_03798_),
    .B1(_05250_),
    .Y(_03864_));
 sky130_fd_sc_hd__a31oi_2 _15693_ (.A1(_03809_),
    .A2(net403),
    .A3(_03787_),
    .B1(_01995_),
    .Y(_03875_));
 sky130_fd_sc_hd__a31o_2 _15694_ (.A1(_03809_),
    .A2(net403),
    .A3(_03787_),
    .B1(_01995_),
    .X(_03886_));
 sky130_fd_sc_hd__a22o_1 _15695_ (.A1(net1),
    .A2(_01897_),
    .B1(_03842_),
    .B2(_03864_),
    .X(_03897_));
 sky130_fd_sc_hd__nand4_2 _15696_ (.A(_03864_),
    .B(net1),
    .C(_03842_),
    .D(_01897_),
    .Y(_03908_));
 sky130_fd_sc_hd__o211ai_4 _15697_ (.A1(net305),
    .A2(net303),
    .B1(_03897_),
    .C1(_03908_),
    .Y(_03919_));
 sky130_fd_sc_hd__or4_4 _15698_ (.A(net305),
    .B(net303),
    .C(_03776_),
    .D(_03798_),
    .X(_03930_));
 sky130_fd_sc_hd__a21oi_2 _15699_ (.A1(_03919_),
    .A2(_03930_),
    .B1(_03289_),
    .Y(_03941_));
 sky130_fd_sc_hd__a21o_2 _15700_ (.A1(_03919_),
    .A2(_03930_),
    .B1(_03289_),
    .X(_03953_));
 sky130_fd_sc_hd__and3_1 _15701_ (.A(_03289_),
    .B(_03919_),
    .C(_03930_),
    .X(_03964_));
 sky130_fd_sc_hd__or4_4 _15702_ (.A(net64),
    .B(net34),
    .C(net35),
    .D(_12659_),
    .X(_03975_));
 sky130_fd_sc_hd__o311a_4 _15703_ (.A1(net34),
    .A2(net35),
    .A3(_14447_),
    .B1(net36),
    .C1(net409),
    .X(_03986_));
 sky130_fd_sc_hd__a21oi_4 _15704_ (.A1(_03975_),
    .A2(net409),
    .B1(net36),
    .Y(_03997_));
 sky130_fd_sc_hd__a21boi_4 _15705_ (.A1(_03975_),
    .A2(net409),
    .B1_N(net36),
    .Y(_04008_));
 sky130_fd_sc_hd__and3b_4 _15706_ (.A_N(net36),
    .B(_03975_),
    .C(net409),
    .X(_04019_));
 sky130_fd_sc_hd__nor2_8 _15707_ (.A(_03986_),
    .B(_03997_),
    .Y(_04029_));
 sky130_fd_sc_hd__nor2_8 _15708_ (.A(_04008_),
    .B(net300),
    .Y(_04040_));
 sky130_fd_sc_hd__o22a_1 _15709_ (.A1(_03941_),
    .A2(_03964_),
    .B1(net301),
    .B2(net300),
    .X(_04051_));
 sky130_fd_sc_hd__a31o_1 _15710_ (.A1(_03919_),
    .A2(_03930_),
    .A3(_04040_),
    .B1(_04051_),
    .X(_04063_));
 sky130_fd_sc_hd__o21ai_1 _15711_ (.A1(_05051_),
    .A2(_02027_),
    .B1(_04063_),
    .Y(_04074_));
 sky130_fd_sc_hd__or3_1 _15712_ (.A(_05051_),
    .B(_02027_),
    .C(_04063_),
    .X(_04085_));
 sky130_fd_sc_hd__and2_1 _15713_ (.A(_04074_),
    .B(_04085_),
    .X(net68));
 sky130_fd_sc_hd__o2bb2a_1 _15714_ (.A1_N(_02027_),
    .A2_N(_04063_),
    .B1(_04832_),
    .B2(_04942_),
    .X(_04106_));
 sky130_fd_sc_hd__a21oi_2 _15715_ (.A1(_03400_),
    .A2(_03388_),
    .B1(_03356_),
    .Y(_04117_));
 sky130_fd_sc_hd__o32ai_4 _15716_ (.A1(net380),
    .A2(net391),
    .A3(_03323_),
    .B1(_03411_),
    .B2(_03378_),
    .Y(_04128_));
 sky130_fd_sc_hd__and3_1 _15717_ (.A(_00152_),
    .B(_04503_),
    .C(_04392_),
    .X(_04139_));
 sky130_fd_sc_hd__or3_2 _15718_ (.A(net3),
    .B(net4),
    .C(_00163_),
    .X(_04150_));
 sky130_fd_sc_hd__a311oi_4 _15719_ (.A1(_00152_),
    .A2(_04503_),
    .A3(_04392_),
    .B1(_03399_),
    .C1(net5),
    .Y(_04161_));
 sky130_fd_sc_hd__a311o_4 _15720_ (.A1(_00152_),
    .A2(_04503_),
    .A3(_04392_),
    .B1(_03399_),
    .C1(net5),
    .X(_04173_));
 sky130_fd_sc_hd__o21a_4 _15721_ (.A1(_03399_),
    .A2(_04139_),
    .B1(net5),
    .X(_04184_));
 sky130_fd_sc_hd__o21ai_4 _15722_ (.A1(_03399_),
    .A2(_04139_),
    .B1(net5),
    .Y(_04195_));
 sky130_fd_sc_hd__o311a_4 _15723_ (.A1(net3),
    .A2(net4),
    .A3(_00163_),
    .B1(net5),
    .C1(net410),
    .X(_04206_));
 sky130_fd_sc_hd__a21oi_4 _15724_ (.A1(_04150_),
    .A2(net410),
    .B1(net5),
    .Y(_04216_));
 sky130_fd_sc_hd__or2_4 _15725_ (.A(_04206_),
    .B(_04216_),
    .X(_04227_));
 sky130_fd_sc_hd__nor2_8 _15726_ (.A(_04206_),
    .B(_04216_),
    .Y(_04238_));
 sky130_fd_sc_hd__or3_4 _15727_ (.A(_03178_),
    .B(_04206_),
    .C(_04216_),
    .X(_04249_));
 sky130_fd_sc_hd__o221a_1 _15728_ (.A1(net408),
    .A2(_05152_),
    .B1(_04161_),
    .B2(_04184_),
    .C1(net33),
    .X(_04260_));
 sky130_fd_sc_hd__or4_2 _15729_ (.A(_03178_),
    .B(_05174_),
    .C(_04206_),
    .D(_04216_),
    .X(_04271_));
 sky130_fd_sc_hd__o32a_1 _15730_ (.A1(_03178_),
    .A2(_04206_),
    .A3(_04216_),
    .B1(_02093_),
    .B2(_02115_),
    .X(_04283_));
 sky130_fd_sc_hd__a22o_1 _15731_ (.A1(_02104_),
    .A2(_02126_),
    .B1(net298),
    .B2(net33),
    .X(_04294_));
 sky130_fd_sc_hd__o221a_2 _15732_ (.A1(_02049_),
    .A2(net342),
    .B1(_04161_),
    .B2(_04184_),
    .C1(net33),
    .X(_04305_));
 sky130_fd_sc_hd__o31a_2 _15733_ (.A1(_04206_),
    .A2(_04216_),
    .A3(_02159_),
    .B1(_04294_),
    .X(_04316_));
 sky130_fd_sc_hd__o21ai_4 _15734_ (.A1(net299),
    .A2(_02159_),
    .B1(_04294_),
    .Y(_04327_));
 sky130_fd_sc_hd__nor4_2 _15735_ (.A(_11397_),
    .B(_12987_),
    .C(_00306_),
    .D(_02214_),
    .Y(_04338_));
 sky130_fd_sc_hd__inv_2 _15736_ (.A(_04338_),
    .Y(_04349_));
 sky130_fd_sc_hd__a21oi_2 _15737_ (.A1(_00262_),
    .A2(_02148_),
    .B1(_04338_),
    .Y(_04360_));
 sky130_fd_sc_hd__nand2_2 _15738_ (.A(_02247_),
    .B(_04360_),
    .Y(_04371_));
 sky130_fd_sc_hd__o21a_1 _15739_ (.A1(_11430_),
    .A2(_11473_),
    .B1(_04338_),
    .X(_04381_));
 sky130_fd_sc_hd__o21ai_2 _15740_ (.A1(_11430_),
    .A2(_11473_),
    .B1(_04338_),
    .Y(_04393_));
 sky130_fd_sc_hd__o2bb2ai_4 _15741_ (.A1_N(_04360_),
    .A2_N(_02247_),
    .B1(_11506_),
    .B2(_04349_),
    .Y(_04404_));
 sky130_fd_sc_hd__o21ai_4 _15742_ (.A1(_04283_),
    .A2(_04305_),
    .B1(_04404_),
    .Y(_04415_));
 sky130_fd_sc_hd__a211oi_2 _15743_ (.A1(_02247_),
    .A2(_04360_),
    .B1(_04381_),
    .C1(_04327_),
    .Y(_04426_));
 sky130_fd_sc_hd__o211ai_4 _15744_ (.A1(_11506_),
    .A2(_04349_),
    .B1(_04316_),
    .C1(_04371_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand2_1 _15745_ (.A(_04415_),
    .B(_04437_),
    .Y(_04448_));
 sky130_fd_sc_hd__nand3_2 _15746_ (.A(_04415_),
    .B(_04437_),
    .C(_05174_),
    .Y(_04459_));
 sky130_fd_sc_hd__o32a_1 _15747_ (.A1(_03178_),
    .A2(_04206_),
    .A3(_04216_),
    .B1(net408),
    .B2(_05152_),
    .X(_04470_));
 sky130_fd_sc_hd__a21oi_4 _15748_ (.A1(_04415_),
    .A2(_04437_),
    .B1(_05185_),
    .Y(_04481_));
 sky130_fd_sc_hd__a31o_1 _15749_ (.A1(_05141_),
    .A2(_05163_),
    .A3(_04448_),
    .B1(_04470_),
    .X(_04492_));
 sky130_fd_sc_hd__a21oi_2 _15750_ (.A1(_04271_),
    .A2(_04459_),
    .B1(net388),
    .Y(_04504_));
 sky130_fd_sc_hd__or4_2 _15751_ (.A(net402),
    .B(net400),
    .C(_04470_),
    .D(_04481_),
    .X(_04515_));
 sky130_fd_sc_hd__a311oi_4 _15752_ (.A1(_04415_),
    .A2(_04437_),
    .A3(_05174_),
    .B1(net319),
    .C1(_04260_),
    .Y(_04526_));
 sky130_fd_sc_hd__nand3_4 _15753_ (.A(_04459_),
    .B(net320),
    .C(_04271_),
    .Y(_04536_));
 sky130_fd_sc_hd__or3_4 _15754_ (.A(_00218_),
    .B(_00229_),
    .C(_04470_),
    .X(_04547_));
 sky130_fd_sc_hd__a21oi_1 _15755_ (.A1(_04448_),
    .A2(_05174_),
    .B1(_04547_),
    .Y(_04558_));
 sky130_fd_sc_hd__a21o_1 _15756_ (.A1(_04448_),
    .A2(_05174_),
    .B1(_04547_),
    .X(_04569_));
 sky130_fd_sc_hd__o21a_1 _15757_ (.A1(_04547_),
    .A2(_04481_),
    .B1(_04536_),
    .X(_04580_));
 sky130_fd_sc_hd__o21ai_4 _15758_ (.A1(_04547_),
    .A2(_04481_),
    .B1(_04536_),
    .Y(_04591_));
 sky130_fd_sc_hd__a22oi_4 _15759_ (.A1(_02290_),
    .A2(_02367_),
    .B1(_02444_),
    .B2(_02356_),
    .Y(_04602_));
 sky130_fd_sc_hd__o22ai_4 _15760_ (.A1(_02378_),
    .A2(_02279_),
    .B1(_02345_),
    .B2(_02433_),
    .Y(_04614_));
 sky130_fd_sc_hd__o211ai_4 _15761_ (.A1(_04547_),
    .A2(_04481_),
    .B1(_04536_),
    .C1(_04614_),
    .Y(_04625_));
 sky130_fd_sc_hd__o21a_1 _15762_ (.A1(_04526_),
    .A2(_04558_),
    .B1(_04602_),
    .X(_04636_));
 sky130_fd_sc_hd__o21ai_1 _15763_ (.A1(_04526_),
    .A2(_04558_),
    .B1(_04602_),
    .Y(_04647_));
 sky130_fd_sc_hd__o22ai_2 _15764_ (.A1(net402),
    .A2(net400),
    .B1(_04602_),
    .B2(_04591_),
    .Y(_04658_));
 sky130_fd_sc_hd__o211ai_2 _15765_ (.A1(net402),
    .A2(net400),
    .B1(_04625_),
    .C1(_04647_),
    .Y(_04668_));
 sky130_fd_sc_hd__o22ai_4 _15766_ (.A1(net388),
    .A2(_04492_),
    .B1(_04636_),
    .B2(_04658_),
    .Y(_04679_));
 sky130_fd_sc_hd__a21oi_2 _15767_ (.A1(_02586_),
    .A2(_02608_),
    .B1(_02532_),
    .Y(_04690_));
 sky130_fd_sc_hd__o21ai_2 _15768_ (.A1(_02575_),
    .A2(_02597_),
    .B1(_02543_),
    .Y(_04701_));
 sky130_fd_sc_hd__o22a_1 _15769_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_04636_),
    .B2(_04658_),
    .X(_04712_));
 sky130_fd_sc_hd__a31o_1 _15770_ (.A1(net388),
    .A2(_04625_),
    .A3(_04647_),
    .B1(net325),
    .X(_04723_));
 sky130_fd_sc_hd__o311a_2 _15771_ (.A1(net388),
    .A2(_04470_),
    .A3(_04481_),
    .B1(_12888_),
    .C1(_04668_),
    .X(_04734_));
 sky130_fd_sc_hd__a21oi_1 _15772_ (.A1(_04515_),
    .A2(_04668_),
    .B1(_12888_),
    .Y(_04745_));
 sky130_fd_sc_hd__o21ai_4 _15773_ (.A1(_12845_),
    .A2(_12856_),
    .B1(_04679_),
    .Y(_04756_));
 sky130_fd_sc_hd__o211ai_4 _15774_ (.A1(_04504_),
    .A2(_04723_),
    .B1(_04756_),
    .C1(_04701_),
    .Y(_04767_));
 sky130_fd_sc_hd__o21ai_2 _15775_ (.A1(_04734_),
    .A2(_04745_),
    .B1(_04690_),
    .Y(_04778_));
 sky130_fd_sc_hd__and3_1 _15776_ (.A(_05687_),
    .B(_05709_),
    .C(_04679_),
    .X(_04788_));
 sky130_fd_sc_hd__a211o_2 _15777_ (.A1(_04515_),
    .A2(_04668_),
    .B1(net384),
    .C1(net383),
    .X(_04799_));
 sky130_fd_sc_hd__o211a_1 _15778_ (.A1(net384),
    .A2(net383),
    .B1(_04767_),
    .C1(_04778_),
    .X(_04810_));
 sky130_fd_sc_hd__nand3_4 _15779_ (.A(_04778_),
    .B(_05720_),
    .C(_04767_),
    .Y(_04821_));
 sky130_fd_sc_hd__a31o_2 _15780_ (.A1(_04778_),
    .A2(_05720_),
    .A3(_04767_),
    .B1(_04788_),
    .X(_04833_));
 sky130_fd_sc_hd__a2bb2oi_4 _15781_ (.A1_N(_11210_),
    .A2_N(_11232_),
    .B1(_04799_),
    .B2(_04821_),
    .Y(_04844_));
 sky130_fd_sc_hd__o22ai_4 _15782_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_04788_),
    .B2(_04810_),
    .Y(_04855_));
 sky130_fd_sc_hd__o211a_2 _15783_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_04799_),
    .C1(_04821_),
    .X(_04866_));
 sky130_fd_sc_hd__o211ai_4 _15784_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_04799_),
    .C1(_04821_),
    .Y(_04877_));
 sky130_fd_sc_hd__o21ai_2 _15785_ (.A1(_02685_),
    .A2(_02718_),
    .B1(_02751_),
    .Y(_04887_));
 sky130_fd_sc_hd__o22a_1 _15786_ (.A1(_02510_),
    .A2(_02729_),
    .B1(_02685_),
    .B2(_02718_),
    .X(_04898_));
 sky130_fd_sc_hd__nand3_2 _15787_ (.A(_04855_),
    .B(_04877_),
    .C(_04898_),
    .Y(_04909_));
 sky130_fd_sc_hd__o21ai_2 _15788_ (.A1(_04844_),
    .A2(_04866_),
    .B1(_04887_),
    .Y(_04920_));
 sky130_fd_sc_hd__nand3_1 _15789_ (.A(_04855_),
    .B(_04877_),
    .C(_04887_),
    .Y(_04931_));
 sky130_fd_sc_hd__o2bb2ai_1 _15790_ (.A1_N(_02696_),
    .A2_N(_02762_),
    .B1(_04844_),
    .B2(_04866_),
    .Y(_04943_));
 sky130_fd_sc_hd__nand3_1 _15791_ (.A(_04943_),
    .B(_06837_),
    .C(_04931_),
    .Y(_04954_));
 sky130_fd_sc_hd__and3_1 _15792_ (.A(_04833_),
    .B(_06826_),
    .C(_06804_),
    .X(_04964_));
 sky130_fd_sc_hd__a211o_1 _15793_ (.A1(_04799_),
    .A2(_04821_),
    .B1(net379),
    .C1(net378),
    .X(_04975_));
 sky130_fd_sc_hd__nand3_1 _15794_ (.A(_04920_),
    .B(_06837_),
    .C(_04909_),
    .Y(_04986_));
 sky130_fd_sc_hd__a31o_2 _15795_ (.A1(_04920_),
    .A2(_06837_),
    .A3(_04909_),
    .B1(_04964_),
    .X(_04997_));
 sky130_fd_sc_hd__a311o_1 _15796_ (.A1(_04909_),
    .A2(_04920_),
    .A3(_06837_),
    .B1(_04964_),
    .C1(net356),
    .X(_05008_));
 sky130_fd_sc_hd__o221ai_4 _15797_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_04833_),
    .B2(_06837_),
    .C1(_04954_),
    .Y(_05019_));
 sky130_fd_sc_hd__a31o_1 _15798_ (.A1(_04920_),
    .A2(_06837_),
    .A3(_04909_),
    .B1(net348),
    .X(_05029_));
 sky130_fd_sc_hd__and3_1 _15799_ (.A(_04986_),
    .B(_10015_),
    .C(_04975_),
    .X(_05040_));
 sky130_fd_sc_hd__nand3_1 _15800_ (.A(_04986_),
    .B(_10015_),
    .C(_04975_),
    .Y(_05052_));
 sky130_fd_sc_hd__a32oi_1 _15801_ (.A1(_08907_),
    .A2(_02806_),
    .A3(_02828_),
    .B1(_00931_),
    .B2(_01052_),
    .Y(_05063_));
 sky130_fd_sc_hd__o22ai_4 _15802_ (.A1(_02817_),
    .A2(_02937_),
    .B1(_02959_),
    .B2(_02871_),
    .Y(_05073_));
 sky130_fd_sc_hd__o2111a_1 _15803_ (.A1(_02860_),
    .A2(_02948_),
    .B1(_02970_),
    .C1(_05019_),
    .D1(_05052_),
    .X(_05084_));
 sky130_fd_sc_hd__o2111ai_1 _15804_ (.A1(_02860_),
    .A2(_02948_),
    .B1(_02970_),
    .C1(_05019_),
    .D1(_05052_),
    .Y(_05095_));
 sky130_fd_sc_hd__a21oi_1 _15805_ (.A1(_05019_),
    .A2(_05052_),
    .B1(_05073_),
    .Y(_05105_));
 sky130_fd_sc_hd__o2bb2ai_1 _15806_ (.A1_N(_05019_),
    .A2_N(_05052_),
    .B1(_05063_),
    .B2(_02959_),
    .Y(_05115_));
 sky130_fd_sc_hd__nand3_2 _15807_ (.A(_05115_),
    .B(_07713_),
    .C(_05095_),
    .Y(_05116_));
 sky130_fd_sc_hd__a211o_1 _15808_ (.A1(_04975_),
    .A2(_04986_),
    .B1(net372),
    .C1(net371),
    .X(_05117_));
 sky130_fd_sc_hd__o22ai_1 _15809_ (.A1(net372),
    .A2(net371),
    .B1(_05084_),
    .B2(_05105_),
    .Y(_05118_));
 sky130_fd_sc_hd__o21ai_4 _15810_ (.A1(_07713_),
    .A2(_04997_),
    .B1(_05116_),
    .Y(_05120_));
 sky130_fd_sc_hd__o311a_1 _15811_ (.A1(_07724_),
    .A2(_05084_),
    .A3(_05105_),
    .B1(_08732_),
    .C1(_05008_),
    .X(_05121_));
 sky130_fd_sc_hd__or3_2 _15812_ (.A(net353),
    .B(net352),
    .C(_05120_),
    .X(_05122_));
 sky130_fd_sc_hd__o311a_1 _15813_ (.A1(_06989_),
    .A2(_07011_),
    .A3(_01140_),
    .B1(_03047_),
    .C1(_03091_),
    .X(_05123_));
 sky130_fd_sc_hd__o211ai_1 _15814_ (.A1(_07033_),
    .A2(_01140_),
    .B1(_03047_),
    .C1(_03091_),
    .Y(_05124_));
 sky130_fd_sc_hd__a31oi_4 _15815_ (.A1(_01206_),
    .A2(_03047_),
    .A3(_03091_),
    .B1(_03058_),
    .Y(_05125_));
 sky130_fd_sc_hd__o21ai_2 _15816_ (.A1(_07899_),
    .A2(_03014_),
    .B1(_05124_),
    .Y(_05126_));
 sky130_fd_sc_hd__a21oi_2 _15817_ (.A1(_05008_),
    .A2(_05116_),
    .B1(_08918_),
    .Y(_05127_));
 sky130_fd_sc_hd__nand3_2 _15818_ (.A(_05118_),
    .B(_08907_),
    .C(_05117_),
    .Y(_05128_));
 sky130_fd_sc_hd__o211a_1 _15819_ (.A1(_07713_),
    .A2(_04997_),
    .B1(_05116_),
    .C1(_08918_),
    .X(_05129_));
 sky130_fd_sc_hd__o211ai_2 _15820_ (.A1(_07713_),
    .A2(_04997_),
    .B1(_05116_),
    .C1(_08918_),
    .Y(_05131_));
 sky130_fd_sc_hd__o22ai_1 _15821_ (.A1(_03080_),
    .A2(_03102_),
    .B1(_05127_),
    .B2(_05129_),
    .Y(_05132_));
 sky130_fd_sc_hd__nand3_1 _15822_ (.A(_05126_),
    .B(_05128_),
    .C(_05131_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand3_2 _15823_ (.A(_05125_),
    .B(_05128_),
    .C(_05131_),
    .Y(_05134_));
 sky130_fd_sc_hd__o22ai_2 _15824_ (.A1(_03058_),
    .A2(_05123_),
    .B1(_05127_),
    .B2(_05129_),
    .Y(_05135_));
 sky130_fd_sc_hd__a22oi_2 _15825_ (.A1(_08689_),
    .A2(_08711_),
    .B1(_05132_),
    .B2(_05133_),
    .Y(_05136_));
 sky130_fd_sc_hd__nand3_4 _15826_ (.A(_05135_),
    .B(_08721_),
    .C(_05134_),
    .Y(_05137_));
 sky130_fd_sc_hd__a31o_1 _15827_ (.A1(_05135_),
    .A2(_08721_),
    .A3(_05134_),
    .B1(_05121_),
    .X(_05138_));
 sky130_fd_sc_hd__and3_1 _15828_ (.A(_09796_),
    .B(_09818_),
    .C(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__a2bb2oi_4 _15829_ (.A1_N(net389),
    .A2_N(net370),
    .B1(_05122_),
    .B2(_05137_),
    .Y(_05140_));
 sky130_fd_sc_hd__o22ai_4 _15830_ (.A1(net389),
    .A2(net370),
    .B1(_05121_),
    .B2(_05136_),
    .Y(_05142_));
 sky130_fd_sc_hd__o221a_2 _15831_ (.A1(net369),
    .A2(_07866_),
    .B1(_08721_),
    .B2(_05120_),
    .C1(_05137_),
    .X(_05143_));
 sky130_fd_sc_hd__nand3_4 _15832_ (.A(_05137_),
    .B(_07888_),
    .C(_05122_),
    .Y(_05144_));
 sky130_fd_sc_hd__o221ai_4 _15833_ (.A1(_06332_),
    .A2(_01293_),
    .B1(_07033_),
    .B2(_03179_),
    .C1(_01403_),
    .Y(_05145_));
 sky130_fd_sc_hd__o32a_1 _15834_ (.A1(_06945_),
    .A2(net377),
    .A3(_03167_),
    .B1(_03256_),
    .B2(_03223_),
    .X(_05146_));
 sky130_fd_sc_hd__a21oi_2 _15835_ (.A1(_03223_),
    .A2(_03245_),
    .B1(_03256_),
    .Y(_05147_));
 sky130_fd_sc_hd__o21ai_4 _15836_ (.A1(_05140_),
    .A2(_05143_),
    .B1(_05146_),
    .Y(_05148_));
 sky130_fd_sc_hd__nand3_4 _15837_ (.A(_05142_),
    .B(_05144_),
    .C(_05147_),
    .Y(_05149_));
 sky130_fd_sc_hd__o21ai_2 _15838_ (.A1(_05140_),
    .A2(_05143_),
    .B1(_05147_),
    .Y(_05150_));
 sky130_fd_sc_hd__o211ai_4 _15839_ (.A1(_03167_),
    .A2(_07044_),
    .B1(_05145_),
    .C1(_05144_),
    .Y(_05151_));
 sky130_fd_sc_hd__nand4_2 _15840_ (.A(_03245_),
    .B(_05142_),
    .C(_05144_),
    .D(_05145_),
    .Y(_05153_));
 sky130_fd_sc_hd__nand3_1 _15841_ (.A(_05150_),
    .B(_05153_),
    .C(net337),
    .Y(_05154_));
 sky130_fd_sc_hd__nand3_2 _15842_ (.A(_05148_),
    .B(_05149_),
    .C(_09829_),
    .Y(_05155_));
 sky130_fd_sc_hd__o311a_2 _15843_ (.A1(net353),
    .A2(_05120_),
    .A3(net352),
    .B1(_09840_),
    .C1(_05137_),
    .X(_05156_));
 sky130_fd_sc_hd__inv_2 _15844_ (.A(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__a31oi_4 _15845_ (.A1(_05150_),
    .A2(_05153_),
    .A3(net337),
    .B1(_05139_),
    .Y(_05158_));
 sky130_fd_sc_hd__a31oi_4 _15846_ (.A1(_05148_),
    .A2(_05149_),
    .A3(_09829_),
    .B1(_05156_),
    .Y(_05159_));
 sky130_fd_sc_hd__a22oi_4 _15847_ (.A1(_07000_),
    .A2(_07022_),
    .B1(_05155_),
    .B2(_05157_),
    .Y(_05160_));
 sky130_fd_sc_hd__nand3b_1 _15848_ (.A_N(_05139_),
    .B(_05154_),
    .C(_07033_),
    .Y(_05161_));
 sky130_fd_sc_hd__a311oi_4 _15849_ (.A1(_05148_),
    .A2(_05149_),
    .A3(_09829_),
    .B1(_05156_),
    .C1(_07033_),
    .Y(_05162_));
 sky130_fd_sc_hd__o211ai_4 _15850_ (.A1(_05138_),
    .A2(net337),
    .B1(_07044_),
    .C1(_05155_),
    .Y(_05164_));
 sky130_fd_sc_hd__and3_1 _15851_ (.A(_04128_),
    .B(_05161_),
    .C(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__nand3_1 _15852_ (.A(_04128_),
    .B(_05161_),
    .C(_05164_),
    .Y(_05166_));
 sky130_fd_sc_hd__o221a_1 _15853_ (.A1(_03411_),
    .A2(_03378_),
    .B1(_05162_),
    .B2(_05160_),
    .C1(_03367_),
    .X(_05167_));
 sky130_fd_sc_hd__a21o_1 _15854_ (.A1(_05161_),
    .A2(_05164_),
    .B1(_04128_),
    .X(_05168_));
 sky130_fd_sc_hd__o22ai_2 _15855_ (.A1(net347),
    .A2(net346),
    .B1(_05165_),
    .B2(_05167_),
    .Y(_05169_));
 sky130_fd_sc_hd__a311o_1 _15856_ (.A1(_05148_),
    .A2(_05149_),
    .A3(_09829_),
    .B1(_05156_),
    .C1(_11068_),
    .X(_05170_));
 sky130_fd_sc_hd__nand3_4 _15857_ (.A(_05168_),
    .B(_11068_),
    .C(_05166_),
    .Y(_05171_));
 sky130_fd_sc_hd__o21ai_2 _15858_ (.A1(_11068_),
    .A2(_05158_),
    .B1(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__a211o_2 _15859_ (.A1(_05170_),
    .A2(_05171_),
    .B1(net328),
    .C1(_12681_),
    .X(_05173_));
 sky130_fd_sc_hd__a2bb2oi_2 _15860_ (.A1_N(net392),
    .A2_N(net382),
    .B1(_05170_),
    .B2(_05171_),
    .Y(_05175_));
 sky130_fd_sc_hd__o221ai_4 _15861_ (.A1(net392),
    .A2(net382),
    .B1(_11068_),
    .B2(_05159_),
    .C1(_05169_),
    .Y(_05176_));
 sky130_fd_sc_hd__o221a_1 _15862_ (.A1(net380),
    .A2(net391),
    .B1(_11068_),
    .B2(_05158_),
    .C1(_05171_),
    .X(_05177_));
 sky130_fd_sc_hd__o221ai_4 _15863_ (.A1(net380),
    .A2(net391),
    .B1(_11068_),
    .B2(_05158_),
    .C1(_05171_),
    .Y(_05178_));
 sky130_fd_sc_hd__a22oi_4 _15864_ (.A1(_03345_),
    .A2(_03643_),
    .B1(_03632_),
    .B2(_03533_),
    .Y(_05179_));
 sky130_fd_sc_hd__a22o_1 _15865_ (.A1(_03345_),
    .A2(_03643_),
    .B1(_03632_),
    .B2(_03533_),
    .X(_05180_));
 sky130_fd_sc_hd__o21ai_1 _15866_ (.A1(_05175_),
    .A2(_05177_),
    .B1(_05179_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand3_1 _15867_ (.A(_05176_),
    .B(_05178_),
    .C(_05180_),
    .Y(_05182_));
 sky130_fd_sc_hd__o21ai_1 _15868_ (.A1(_05175_),
    .A2(_05177_),
    .B1(_05180_),
    .Y(_05183_));
 sky130_fd_sc_hd__nand2_1 _15869_ (.A(_05179_),
    .B(_05178_),
    .Y(_05184_));
 sky130_fd_sc_hd__o211ai_2 _15870_ (.A1(_06343_),
    .A2(_05172_),
    .B1(_05179_),
    .C1(_05176_),
    .Y(_05186_));
 sky130_fd_sc_hd__nand3_1 _15871_ (.A(_05181_),
    .B(_05182_),
    .C(net313),
    .Y(_05187_));
 sky130_fd_sc_hd__o311a_1 _15872_ (.A1(_11079_),
    .A2(_05165_),
    .A3(_05167_),
    .B1(_05170_),
    .C1(_12703_),
    .X(_05188_));
 sky130_fd_sc_hd__a31o_1 _15873_ (.A1(_05181_),
    .A2(_05182_),
    .A3(net313),
    .B1(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__o31a_2 _15874_ (.A1(net328),
    .A2(_12681_),
    .A3(_05172_),
    .B1(_05187_),
    .X(_05190_));
 sky130_fd_sc_hd__a31oi_2 _15875_ (.A1(_01853_),
    .A2(net386),
    .A3(_01798_),
    .B1(_03709_),
    .Y(_05191_));
 sky130_fd_sc_hd__a32oi_4 _15876_ (.A1(_03698_),
    .A2(_05534_),
    .A3(_05512_),
    .B1(_03820_),
    .B2(_03732_),
    .Y(_05192_));
 sky130_fd_sc_hd__o211ai_4 _15877_ (.A1(_03709_),
    .A2(_03720_),
    .B1(_03765_),
    .C1(_03831_),
    .Y(_05193_));
 sky130_fd_sc_hd__o2111a_1 _15878_ (.A1(_03709_),
    .A2(_03720_),
    .B1(_03831_),
    .C1(_05851_),
    .D1(_03765_),
    .X(_05194_));
 sky130_fd_sc_hd__o2111ai_4 _15879_ (.A1(_03709_),
    .A2(_03720_),
    .B1(_03831_),
    .C1(_05851_),
    .D1(_03765_),
    .Y(_05195_));
 sky130_fd_sc_hd__o22a_1 _15880_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_03754_),
    .B2(_05191_),
    .X(_05197_));
 sky130_fd_sc_hd__o22ai_4 _15881_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_03754_),
    .B2(_05191_),
    .Y(_05198_));
 sky130_fd_sc_hd__a31oi_2 _15882_ (.A1(_05198_),
    .A2(_00055_),
    .A3(_05195_),
    .B1(_05190_),
    .Y(_05199_));
 sky130_fd_sc_hd__a31o_1 _15883_ (.A1(_05198_),
    .A2(_00055_),
    .A3(_05195_),
    .B1(_05190_),
    .X(_05200_));
 sky130_fd_sc_hd__nand4_1 _15884_ (.A(_05190_),
    .B(_05195_),
    .C(_05198_),
    .D(_00055_),
    .Y(_05201_));
 sky130_fd_sc_hd__a31oi_4 _15885_ (.A1(_05183_),
    .A2(_05186_),
    .A3(net313),
    .B1(_05862_),
    .Y(_05202_));
 sky130_fd_sc_hd__a311oi_2 _15886_ (.A1(_05181_),
    .A2(_05182_),
    .A3(net313),
    .B1(_05188_),
    .C1(_05851_),
    .Y(_05203_));
 sky130_fd_sc_hd__o211ai_2 _15887_ (.A1(net313),
    .A2(_05172_),
    .B1(_05187_),
    .C1(_05862_),
    .Y(_05204_));
 sky130_fd_sc_hd__a41oi_4 _15888_ (.A1(_00055_),
    .A2(_05190_),
    .A3(_05195_),
    .A4(_05198_),
    .B1(_05199_),
    .Y(_05205_));
 sky130_fd_sc_hd__o41ai_2 _15889_ (.A1(_00066_),
    .A2(_05189_),
    .A3(_05194_),
    .A4(_05197_),
    .B1(_05200_),
    .Y(_05206_));
 sky130_fd_sc_hd__o22ai_4 _15890_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_03853_),
    .B2(_03875_),
    .Y(_05208_));
 sky130_fd_sc_hd__o211ai_4 _15891_ (.A1(net398),
    .A2(net397),
    .B1(_03864_),
    .C1(_03886_),
    .Y(_05209_));
 sky130_fd_sc_hd__o2111a_2 _15892_ (.A1(net305),
    .A2(net303),
    .B1(_05209_),
    .C1(_05205_),
    .D1(_05208_),
    .X(_05210_));
 sky130_fd_sc_hd__o2111ai_4 _15893_ (.A1(net305),
    .A2(net303),
    .B1(_05209_),
    .C1(_05205_),
    .D1(_05208_),
    .Y(_05211_));
 sky130_fd_sc_hd__a31oi_4 _15894_ (.A1(_05208_),
    .A2(_05209_),
    .A3(_01962_),
    .B1(_05205_),
    .Y(_05212_));
 sky130_fd_sc_hd__a31o_2 _15895_ (.A1(_05208_),
    .A2(_05209_),
    .A3(_01962_),
    .B1(_05205_),
    .X(_05213_));
 sky130_fd_sc_hd__o2111ai_1 _15896_ (.A1(_03399_),
    .A2(_05491_),
    .B1(_05534_),
    .C1(_05200_),
    .D1(_05201_),
    .Y(_05214_));
 sky130_fd_sc_hd__a21oi_1 _15897_ (.A1(_05211_),
    .A2(_05213_),
    .B1(net275),
    .Y(_05215_));
 sky130_fd_sc_hd__and3_1 _15898_ (.A(_05213_),
    .B(net403),
    .C(_05211_),
    .X(_05216_));
 sky130_fd_sc_hd__nand4_4 _15899_ (.A(_05207_),
    .B(_05229_),
    .C(_05211_),
    .D(_05213_),
    .Y(_05217_));
 sky130_fd_sc_hd__a21oi_2 _15900_ (.A1(_05211_),
    .A2(_05213_),
    .B1(net403),
    .Y(_05219_));
 sky130_fd_sc_hd__o21ai_4 _15901_ (.A1(_05210_),
    .A2(_05212_),
    .B1(_05250_),
    .Y(_05220_));
 sky130_fd_sc_hd__nand3_1 _15902_ (.A(_03953_),
    .B(_05217_),
    .C(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__a221o_1 _15903_ (.A1(_03919_),
    .A2(_03930_),
    .B1(_05217_),
    .B2(_05220_),
    .C1(_03289_),
    .X(_05222_));
 sky130_fd_sc_hd__nand2_2 _15904_ (.A(_05220_),
    .B(_03941_),
    .Y(_05223_));
 sky130_fd_sc_hd__a31oi_2 _15905_ (.A1(_05222_),
    .A2(net275),
    .A3(_05221_),
    .B1(_05215_),
    .Y(_05224_));
 sky130_fd_sc_hd__a311o_4 _15906_ (.A1(_05222_),
    .A2(net275),
    .A3(_05221_),
    .B1(_05215_),
    .C1(_03289_),
    .X(_05225_));
 sky130_fd_sc_hd__nor2_1 _15907_ (.A(net1),
    .B(_05224_),
    .Y(_05226_));
 sky130_fd_sc_hd__or4_4 _15908_ (.A(net34),
    .B(net35),
    .C(net36),
    .D(_14447_),
    .X(_05227_));
 sky130_fd_sc_hd__o311a_4 _15909_ (.A1(net35),
    .A2(net36),
    .A3(_01908_),
    .B1(net37),
    .C1(net409),
    .X(_05228_));
 sky130_fd_sc_hd__a21oi_4 _15910_ (.A1(_05227_),
    .A2(net409),
    .B1(net37),
    .Y(_05230_));
 sky130_fd_sc_hd__a21boi_4 _15911_ (.A1(_05227_),
    .A2(net409),
    .B1_N(net37),
    .Y(_05231_));
 sky130_fd_sc_hd__and3b_4 _15912_ (.A_N(net37),
    .B(_05227_),
    .C(net409),
    .X(_05232_));
 sky130_fd_sc_hd__nor2_8 _15913_ (.A(_05228_),
    .B(_05230_),
    .Y(_05233_));
 sky130_fd_sc_hd__nor2_8 _15914_ (.A(net296),
    .B(_05232_),
    .Y(_05234_));
 sky130_fd_sc_hd__nor3b_1 _15915_ (.A(_05234_),
    .B(_05226_),
    .C_N(_05225_),
    .Y(_05235_));
 sky130_fd_sc_hd__a21oi_1 _15916_ (.A1(_05224_),
    .A2(_05234_),
    .B1(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__xnor2_1 _15917_ (.A(_04106_),
    .B(_05236_),
    .Y(net69));
 sky130_fd_sc_hd__and3_1 _15918_ (.A(_02027_),
    .B(_04063_),
    .C(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__a21oi_4 _15919_ (.A1(_05179_),
    .A2(_05178_),
    .B1(_05175_),
    .Y(_05238_));
 sky130_fd_sc_hd__a21o_1 _15920_ (.A1(_05179_),
    .A2(_05178_),
    .B1(_05175_),
    .X(_05240_));
 sky130_fd_sc_hd__or4_4 _15921_ (.A(net3),
    .B(net4),
    .C(net5),
    .D(_00163_),
    .X(_05241_));
 sky130_fd_sc_hd__and3b_4 _15922_ (.A_N(net6),
    .B(_05241_),
    .C(net410),
    .X(_05242_));
 sky130_fd_sc_hd__or3b_4 _15923_ (.A(_03399_),
    .B(net6),
    .C_N(_05241_),
    .X(_05243_));
 sky130_fd_sc_hd__a21boi_4 _15924_ (.A1(_05241_),
    .A2(net410),
    .B1_N(net6),
    .Y(_05244_));
 sky130_fd_sc_hd__a21bo_4 _15925_ (.A1(_05241_),
    .A2(net410),
    .B1_N(net6),
    .X(_05245_));
 sky130_fd_sc_hd__o311a_4 _15926_ (.A1(net4),
    .A2(net5),
    .A3(_02038_),
    .B1(net6),
    .C1(net410),
    .X(_05246_));
 sky130_fd_sc_hd__a21oi_4 _15927_ (.A1(_05241_),
    .A2(net410),
    .B1(net6),
    .Y(_05247_));
 sky130_fd_sc_hd__nor2_8 _15928_ (.A(net318),
    .B(net315),
    .Y(_05248_));
 sky130_fd_sc_hd__nor2_8 _15929_ (.A(_05246_),
    .B(_05247_),
    .Y(_05249_));
 sky130_fd_sc_hd__o21a_1 _15930_ (.A1(_05242_),
    .A2(net317),
    .B1(net33),
    .X(_05251_));
 sky130_fd_sc_hd__or3_2 _15931_ (.A(_03178_),
    .B(_05246_),
    .C(_05247_),
    .X(_05252_));
 sky130_fd_sc_hd__o221a_2 _15932_ (.A1(net408),
    .A2(_05152_),
    .B1(_05242_),
    .B2(net317),
    .C1(net33),
    .X(_05253_));
 sky130_fd_sc_hd__a31oi_4 _15933_ (.A1(_04371_),
    .A2(_04393_),
    .A3(_04316_),
    .B1(_04305_),
    .Y(_05254_));
 sky130_fd_sc_hd__or3_1 _15934_ (.A(_04161_),
    .B(_04184_),
    .C(_05251_),
    .X(_05255_));
 sky130_fd_sc_hd__or4_1 _15935_ (.A(_03178_),
    .B(_04206_),
    .C(_04216_),
    .D(net295),
    .X(_05256_));
 sky130_fd_sc_hd__o21ai_4 _15936_ (.A1(_04249_),
    .A2(net295),
    .B1(_05255_),
    .Y(_05257_));
 sky130_fd_sc_hd__o21bai_4 _15937_ (.A1(_04305_),
    .A2(_04426_),
    .B1_N(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__o221ai_4 _15938_ (.A1(_02159_),
    .A2(net299),
    .B1(_04327_),
    .B2(_04404_),
    .C1(_05257_),
    .Y(_05259_));
 sky130_fd_sc_hd__o32a_1 _15939_ (.A1(_03178_),
    .A2(_05246_),
    .A3(_05247_),
    .B1(net408),
    .B2(_05152_),
    .X(_05260_));
 sky130_fd_sc_hd__a21oi_1 _15940_ (.A1(_05258_),
    .A2(_05259_),
    .B1(_05185_),
    .Y(_05262_));
 sky130_fd_sc_hd__a21o_1 _15941_ (.A1(_05258_),
    .A2(_05259_),
    .B1(_05185_),
    .X(_05263_));
 sky130_fd_sc_hd__a31oi_4 _15942_ (.A1(_05258_),
    .A2(_05259_),
    .A3(_05174_),
    .B1(_05253_),
    .Y(_05264_));
 sky130_fd_sc_hd__or4_4 _15943_ (.A(net402),
    .B(net400),
    .C(_05260_),
    .D(_05262_),
    .X(_05265_));
 sky130_fd_sc_hd__o22a_1 _15944_ (.A1(_02049_),
    .A2(net342),
    .B1(_05251_),
    .B2(_05174_),
    .X(_05266_));
 sky130_fd_sc_hd__o221a_2 _15945_ (.A1(_02049_),
    .A2(net342),
    .B1(_05251_),
    .B2(_05174_),
    .C1(_05263_),
    .X(_05267_));
 sky130_fd_sc_hd__or4_1 _15946_ (.A(_02093_),
    .B(_02115_),
    .C(_05260_),
    .D(_05262_),
    .X(_05268_));
 sky130_fd_sc_hd__a311oi_4 _15947_ (.A1(_05258_),
    .A2(_05259_),
    .A3(_05174_),
    .B1(_02148_),
    .C1(_05253_),
    .Y(_05269_));
 sky130_fd_sc_hd__a21oi_4 _15948_ (.A1(_05263_),
    .A2(_05266_),
    .B1(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__nand4_2 _15949_ (.A(_02400_),
    .B(_00471_),
    .C(_13229_),
    .D(_02356_),
    .Y(_05271_));
 sky130_fd_sc_hd__nand4_2 _15950_ (.A(_04536_),
    .B(_02411_),
    .C(_00471_),
    .D(_13229_),
    .Y(_05273_));
 sky130_fd_sc_hd__and4b_1 _15951_ (.A_N(_13273_),
    .B(_02400_),
    .C(_00471_),
    .D(_02356_),
    .X(_05274_));
 sky130_fd_sc_hd__nand4b_4 _15952_ (.A_N(_13273_),
    .B(_02400_),
    .C(_00471_),
    .D(_02356_),
    .Y(_05275_));
 sky130_fd_sc_hd__nor3_2 _15953_ (.A(_04526_),
    .B(_05275_),
    .C(_04558_),
    .Y(_05276_));
 sky130_fd_sc_hd__o32a_1 _15954_ (.A1(net320),
    .A2(_04470_),
    .A3(_04481_),
    .B1(_05271_),
    .B2(_04526_),
    .X(_05277_));
 sky130_fd_sc_hd__o22ai_1 _15955_ (.A1(_04481_),
    .A2(_04547_),
    .B1(_05271_),
    .B2(_04526_),
    .Y(_05278_));
 sky130_fd_sc_hd__a21oi_2 _15956_ (.A1(_04580_),
    .A2(_04614_),
    .B1(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__o211ai_4 _15957_ (.A1(_04526_),
    .A2(_04602_),
    .B1(_05273_),
    .C1(_04569_),
    .Y(_05280_));
 sky130_fd_sc_hd__a21oi_4 _15958_ (.A1(_05277_),
    .A2(_04625_),
    .B1(_05276_),
    .Y(_05281_));
 sky130_fd_sc_hd__o311a_1 _15959_ (.A1(_13174_),
    .A2(_04591_),
    .A3(_05271_),
    .B1(_05270_),
    .C1(_05280_),
    .X(_05282_));
 sky130_fd_sc_hd__o211ai_4 _15960_ (.A1(_04591_),
    .A2(_05275_),
    .B1(_05270_),
    .C1(_05280_),
    .Y(_05284_));
 sky130_fd_sc_hd__o22ai_4 _15961_ (.A1(_05267_),
    .A2(_05269_),
    .B1(_05276_),
    .B2(_05279_),
    .Y(_05285_));
 sky130_fd_sc_hd__o22ai_2 _15962_ (.A1(net402),
    .A2(net400),
    .B1(_05270_),
    .B2(_05281_),
    .Y(_05286_));
 sky130_fd_sc_hd__o211ai_4 _15963_ (.A1(net402),
    .A2(net400),
    .B1(_05284_),
    .C1(_05285_),
    .Y(_05287_));
 sky130_fd_sc_hd__o22ai_4 _15964_ (.A1(net388),
    .A2(_05264_),
    .B1(_05282_),
    .B2(_05286_),
    .Y(_05288_));
 sky130_fd_sc_hd__and3_1 _15965_ (.A(_05687_),
    .B(_05709_),
    .C(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__a211o_2 _15966_ (.A1(_05265_),
    .A2(_05287_),
    .B1(net384),
    .C1(net383),
    .X(_05290_));
 sky130_fd_sc_hd__a221oi_4 _15967_ (.A1(_02586_),
    .A2(_02608_),
    .B1(_04679_),
    .B2(net325),
    .C1(_02532_),
    .Y(_05291_));
 sky130_fd_sc_hd__a22oi_4 _15968_ (.A1(_04515_),
    .A2(_04712_),
    .B1(_04690_),
    .B2(_04756_),
    .Y(_05292_));
 sky130_fd_sc_hd__o22ai_2 _15969_ (.A1(_04504_),
    .A2(_04723_),
    .B1(_04745_),
    .B2(_04701_),
    .Y(_05293_));
 sky130_fd_sc_hd__a31oi_2 _15970_ (.A1(net388),
    .A2(_05284_),
    .A3(_05285_),
    .B1(net319),
    .Y(_05295_));
 sky130_fd_sc_hd__o311a_1 _15971_ (.A1(net388),
    .A2(_05260_),
    .A3(_05262_),
    .B1(net320),
    .C1(_05287_),
    .X(_05296_));
 sky130_fd_sc_hd__o211ai_4 _15972_ (.A1(net388),
    .A2(_05264_),
    .B1(net320),
    .C1(_05287_),
    .Y(_05297_));
 sky130_fd_sc_hd__a2bb2oi_4 _15973_ (.A1_N(_00174_),
    .A2_N(_00196_),
    .B1(_05265_),
    .B2(_05287_),
    .Y(_05298_));
 sky130_fd_sc_hd__o21ai_2 _15974_ (.A1(_00174_),
    .A2(_00196_),
    .B1(_05288_),
    .Y(_05299_));
 sky130_fd_sc_hd__a211oi_1 _15975_ (.A1(_05295_),
    .A2(_05265_),
    .B1(_05293_),
    .C1(_05298_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand3_2 _15976_ (.A(_05299_),
    .B(_05292_),
    .C(_05297_),
    .Y(_05301_));
 sky130_fd_sc_hd__a2bb2oi_1 _15977_ (.A1_N(_04734_),
    .A2_N(_05291_),
    .B1(_05297_),
    .B2(_05299_),
    .Y(_05302_));
 sky130_fd_sc_hd__o22ai_4 _15978_ (.A1(_04734_),
    .A2(_05291_),
    .B1(_05296_),
    .B2(_05298_),
    .Y(_05303_));
 sky130_fd_sc_hd__nand3_2 _15979_ (.A(_05303_),
    .B(_05720_),
    .C(_05301_),
    .Y(_05304_));
 sky130_fd_sc_hd__o22ai_2 _15980_ (.A1(net384),
    .A2(net383),
    .B1(_05300_),
    .B2(_05302_),
    .Y(_05306_));
 sky130_fd_sc_hd__a31o_2 _15981_ (.A1(_05303_),
    .A2(_05720_),
    .A3(_05301_),
    .B1(_05289_),
    .X(_05307_));
 sky130_fd_sc_hd__o311a_1 _15982_ (.A1(_05731_),
    .A2(_05300_),
    .A3(_05302_),
    .B1(_06848_),
    .C1(_05290_),
    .X(_05308_));
 sky130_fd_sc_hd__a21oi_2 _15983_ (.A1(net330),
    .A2(_04833_),
    .B1(_04898_),
    .Y(_05309_));
 sky130_fd_sc_hd__o211a_1 _15984_ (.A1(_02685_),
    .A2(_02718_),
    .B1(_02751_),
    .C1(_04877_),
    .X(_05310_));
 sky130_fd_sc_hd__o21ai_1 _15985_ (.A1(_04866_),
    .A2(_04887_),
    .B1(_04855_),
    .Y(_05311_));
 sky130_fd_sc_hd__a311oi_4 _15986_ (.A1(_05303_),
    .A2(_05720_),
    .A3(_05301_),
    .B1(net325),
    .C1(_05289_),
    .Y(_05312_));
 sky130_fd_sc_hd__nand3_4 _15987_ (.A(_05304_),
    .B(_12888_),
    .C(_05290_),
    .Y(_05313_));
 sky130_fd_sc_hd__a2bb2oi_4 _15988_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_05290_),
    .B2(_05304_),
    .Y(_05314_));
 sky130_fd_sc_hd__o211ai_4 _15989_ (.A1(_05288_),
    .A2(net359),
    .B1(net325),
    .C1(_05306_),
    .Y(_05315_));
 sky130_fd_sc_hd__o211ai_4 _15990_ (.A1(_04866_),
    .A2(_05309_),
    .B1(_05313_),
    .C1(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__o22ai_4 _15991_ (.A1(_04844_),
    .A2(_05310_),
    .B1(_05312_),
    .B2(_05314_),
    .Y(_05317_));
 sky130_fd_sc_hd__nand3_2 _15992_ (.A(_05317_),
    .B(net357),
    .C(_05316_),
    .Y(_05318_));
 sky130_fd_sc_hd__o311a_1 _15993_ (.A1(net384),
    .A2(_05288_),
    .A3(net383),
    .B1(_06848_),
    .C1(_05306_),
    .X(_05319_));
 sky130_fd_sc_hd__a211o_1 _15994_ (.A1(_05290_),
    .A2(_05304_),
    .B1(net379),
    .C1(net378),
    .X(_05320_));
 sky130_fd_sc_hd__o211ai_2 _15995_ (.A1(_04844_),
    .A2(_05310_),
    .B1(_05313_),
    .C1(_05315_),
    .Y(_05321_));
 sky130_fd_sc_hd__o22ai_2 _15996_ (.A1(_04866_),
    .A2(_05309_),
    .B1(_05312_),
    .B2(_05314_),
    .Y(_05322_));
 sky130_fd_sc_hd__nand3_1 _15997_ (.A(_05322_),
    .B(net357),
    .C(_05321_),
    .Y(_05323_));
 sky130_fd_sc_hd__a31oi_4 _15998_ (.A1(_05317_),
    .A2(net357),
    .A3(_05316_),
    .B1(_05308_),
    .Y(_05324_));
 sky130_fd_sc_hd__a31oi_4 _15999_ (.A1(_05322_),
    .A2(_06837_),
    .A3(_05321_),
    .B1(_05319_),
    .Y(_05325_));
 sky130_fd_sc_hd__o211a_1 _16000_ (.A1(_05307_),
    .A2(net357),
    .B1(net330),
    .C1(_05318_),
    .X(_05327_));
 sky130_fd_sc_hd__o211ai_4 _16001_ (.A1(_05307_),
    .A2(net357),
    .B1(net330),
    .C1(_05318_),
    .Y(_05328_));
 sky130_fd_sc_hd__and3_1 _16002_ (.A(_05323_),
    .B(net331),
    .C(_05320_),
    .X(_05329_));
 sky130_fd_sc_hd__o211ai_4 _16003_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_05320_),
    .C1(_05323_),
    .Y(_05330_));
 sky130_fd_sc_hd__o211a_1 _16004_ (.A1(_02860_),
    .A2(_02948_),
    .B1(_02970_),
    .C1(_05019_),
    .X(_05331_));
 sky130_fd_sc_hd__a2bb2oi_2 _16005_ (.A1_N(_04964_),
    .A2_N(_05029_),
    .B1(_05073_),
    .B2(_05019_),
    .Y(_05332_));
 sky130_fd_sc_hd__o2bb2ai_1 _16006_ (.A1_N(_05019_),
    .A2_N(_05073_),
    .B1(_05029_),
    .B2(_04964_),
    .Y(_05333_));
 sky130_fd_sc_hd__o211a_4 _16007_ (.A1(_05307_),
    .A2(net357),
    .B1(_07724_),
    .C1(_05318_),
    .X(_05334_));
 sky130_fd_sc_hd__a311o_1 _16008_ (.A1(_05317_),
    .A2(net357),
    .A3(_05316_),
    .B1(net356),
    .C1(_05308_),
    .X(_05335_));
 sky130_fd_sc_hd__a21oi_1 _16009_ (.A1(_05328_),
    .A2(_05330_),
    .B1(_05332_),
    .Y(_05336_));
 sky130_fd_sc_hd__o2bb2ai_2 _16010_ (.A1_N(_05328_),
    .A2_N(_05330_),
    .B1(_05331_),
    .B2(_05040_),
    .Y(_05338_));
 sky130_fd_sc_hd__nand3_2 _16011_ (.A(_05328_),
    .B(_05332_),
    .C(_05330_),
    .Y(_05339_));
 sky130_fd_sc_hd__a31o_1 _16012_ (.A1(_05328_),
    .A2(_05332_),
    .A3(_05330_),
    .B1(_07724_),
    .X(_05340_));
 sky130_fd_sc_hd__nand3_1 _16013_ (.A(_05338_),
    .B(_05339_),
    .C(net356),
    .Y(_05341_));
 sky130_fd_sc_hd__o22ai_4 _16014_ (.A1(net356),
    .A2(_05325_),
    .B1(_05336_),
    .B2(_05340_),
    .Y(_05342_));
 sky130_fd_sc_hd__o311a_2 _16015_ (.A1(net372),
    .A2(_05325_),
    .A3(net371),
    .B1(_08732_),
    .C1(_05341_),
    .X(_05343_));
 sky130_fd_sc_hd__inv_2 _16016_ (.A(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__a2bb2oi_2 _16017_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_05335_),
    .B2(_05341_),
    .Y(_05345_));
 sky130_fd_sc_hd__o21ai_4 _16018_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_05342_),
    .Y(_05346_));
 sky130_fd_sc_hd__a31o_2 _16019_ (.A1(_05338_),
    .A2(_05339_),
    .A3(net356),
    .B1(net348),
    .X(_05347_));
 sky130_fd_sc_hd__a311oi_4 _16020_ (.A1(_05338_),
    .A2(_05339_),
    .A3(net356),
    .B1(net348),
    .C1(_05334_),
    .Y(_05349_));
 sky130_fd_sc_hd__a21oi_4 _16021_ (.A1(_05125_),
    .A2(_05128_),
    .B1(_05129_),
    .Y(_05350_));
 sky130_fd_sc_hd__o32ai_4 _16022_ (.A1(_08863_),
    .A2(net366),
    .A3(_05120_),
    .B1(_05127_),
    .B2(_05126_),
    .Y(_05351_));
 sky130_fd_sc_hd__o21ai_2 _16023_ (.A1(_05345_),
    .A2(_05349_),
    .B1(_05351_),
    .Y(_05352_));
 sky130_fd_sc_hd__o211ai_4 _16024_ (.A1(_05334_),
    .A2(_05347_),
    .B1(_05350_),
    .C1(_05346_),
    .Y(_05353_));
 sky130_fd_sc_hd__and3_1 _16025_ (.A(_05352_),
    .B(_05353_),
    .C(_08721_),
    .X(_05354_));
 sky130_fd_sc_hd__nand3_2 _16026_ (.A(_05352_),
    .B(_05353_),
    .C(_08721_),
    .Y(_05355_));
 sky130_fd_sc_hd__a211o_2 _16027_ (.A1(_05335_),
    .A2(_05341_),
    .B1(net353),
    .C1(net352),
    .X(_05356_));
 sky130_fd_sc_hd__o21ai_1 _16028_ (.A1(_05345_),
    .A2(_05349_),
    .B1(_05350_),
    .Y(_05357_));
 sky130_fd_sc_hd__o211ai_1 _16029_ (.A1(_05334_),
    .A2(_05347_),
    .B1(_05351_),
    .C1(_05346_),
    .Y(_05358_));
 sky130_fd_sc_hd__nand3_2 _16030_ (.A(_05357_),
    .B(_05358_),
    .C(_08721_),
    .Y(_05360_));
 sky130_fd_sc_hd__a31oi_1 _16031_ (.A1(_05352_),
    .A2(_05353_),
    .A3(_08721_),
    .B1(_05343_),
    .Y(_05361_));
 sky130_fd_sc_hd__a31o_1 _16032_ (.A1(_05352_),
    .A2(_05353_),
    .A3(_08721_),
    .B1(_05343_),
    .X(_05362_));
 sky130_fd_sc_hd__a31oi_2 _16033_ (.A1(_03245_),
    .A2(_05144_),
    .A3(_05145_),
    .B1(_05140_),
    .Y(_05363_));
 sky130_fd_sc_hd__a31o_1 _16034_ (.A1(_03245_),
    .A2(_05144_),
    .A3(_05145_),
    .B1(_05140_),
    .X(_05364_));
 sky130_fd_sc_hd__a21oi_1 _16035_ (.A1(_05142_),
    .A2(_05151_),
    .B1(_08907_),
    .Y(_05365_));
 sky130_fd_sc_hd__a31oi_2 _16036_ (.A1(_05151_),
    .A2(_08907_),
    .A3(_05142_),
    .B1(_09840_),
    .Y(_05366_));
 sky130_fd_sc_hd__a31o_1 _16037_ (.A1(_05151_),
    .A2(_08907_),
    .A3(_05142_),
    .B1(_09840_),
    .X(_05367_));
 sky130_fd_sc_hd__o2111ai_4 _16038_ (.A1(_08907_),
    .A2(_05363_),
    .B1(_05355_),
    .C1(_05344_),
    .D1(_05366_),
    .Y(_05368_));
 sky130_fd_sc_hd__o22ai_4 _16039_ (.A1(_05343_),
    .A2(_05354_),
    .B1(_05365_),
    .B2(_05367_),
    .Y(_05369_));
 sky130_fd_sc_hd__o211ai_2 _16040_ (.A1(_08863_),
    .A2(net366),
    .B1(_05356_),
    .C1(_05360_),
    .Y(_05371_));
 sky130_fd_sc_hd__o211a_1 _16041_ (.A1(_08819_),
    .A2(net367),
    .B1(_05344_),
    .C1(_05355_),
    .X(_05372_));
 sky130_fd_sc_hd__o211ai_1 _16042_ (.A1(_08819_),
    .A2(net367),
    .B1(_05344_),
    .C1(_05355_),
    .Y(_05373_));
 sky130_fd_sc_hd__nand3_1 _16043_ (.A(_05364_),
    .B(_05371_),
    .C(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__a21o_1 _16044_ (.A1(_05371_),
    .A2(_05373_),
    .B1(_05364_),
    .X(_05375_));
 sky130_fd_sc_hd__nand3_1 _16045_ (.A(_05375_),
    .B(net337),
    .C(_05374_),
    .Y(_05376_));
 sky130_fd_sc_hd__a311o_2 _16046_ (.A1(_05352_),
    .A2(_05353_),
    .A3(_08721_),
    .B1(net337),
    .C1(_05343_),
    .X(_05377_));
 sky130_fd_sc_hd__and3_4 _16047_ (.A(_11079_),
    .B(_05368_),
    .C(_05369_),
    .X(_05378_));
 sky130_fd_sc_hd__inv_2 _16048_ (.A(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__o211a_1 _16049_ (.A1(_03411_),
    .A2(_03378_),
    .B1(_03367_),
    .C1(_05164_),
    .X(_05380_));
 sky130_fd_sc_hd__a32oi_4 _16050_ (.A1(_06956_),
    .A2(_05158_),
    .A3(_06978_),
    .B1(_04117_),
    .B2(_05164_),
    .Y(_05382_));
 sky130_fd_sc_hd__o32ai_4 _16051_ (.A1(_06945_),
    .A2(net377),
    .A3(_05159_),
    .B1(_05162_),
    .B2(_04128_),
    .Y(_05383_));
 sky130_fd_sc_hd__a31oi_2 _16052_ (.A1(_05375_),
    .A2(net337),
    .A3(_05374_),
    .B1(_07899_),
    .Y(_05384_));
 sky130_fd_sc_hd__a21oi_2 _16053_ (.A1(_05368_),
    .A2(_05369_),
    .B1(_07899_),
    .Y(_05385_));
 sky130_fd_sc_hd__nand3_1 _16054_ (.A(_05376_),
    .B(_05377_),
    .C(_07888_),
    .Y(_05386_));
 sky130_fd_sc_hd__a22oi_2 _16055_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_05376_),
    .B2(_05377_),
    .Y(_05387_));
 sky130_fd_sc_hd__nand3_4 _16056_ (.A(_07899_),
    .B(_05368_),
    .C(_05369_),
    .Y(_05388_));
 sky130_fd_sc_hd__nand3_4 _16057_ (.A(_05382_),
    .B(_05386_),
    .C(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__o22ai_4 _16058_ (.A1(_05160_),
    .A2(_05380_),
    .B1(_05385_),
    .B2(_05387_),
    .Y(_05390_));
 sky130_fd_sc_hd__o211a_1 _16059_ (.A1(net347),
    .A2(net346),
    .B1(_05389_),
    .C1(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__o211ai_4 _16060_ (.A1(net347),
    .A2(net346),
    .B1(_05389_),
    .C1(_05390_),
    .Y(_05393_));
 sky130_fd_sc_hd__a31oi_4 _16061_ (.A1(_05390_),
    .A2(net334),
    .A3(_05389_),
    .B1(_05378_),
    .Y(_05394_));
 sky130_fd_sc_hd__a31o_1 _16062_ (.A1(_05390_),
    .A2(net334),
    .A3(_05389_),
    .B1(_07044_),
    .X(_05395_));
 sky130_fd_sc_hd__a311oi_4 _16063_ (.A1(_05390_),
    .A2(net334),
    .A3(_05389_),
    .B1(_05378_),
    .C1(_07044_),
    .Y(_05396_));
 sky130_fd_sc_hd__a311o_1 _16064_ (.A1(_05390_),
    .A2(net334),
    .A3(_05389_),
    .B1(_05378_),
    .C1(_07044_),
    .X(_05397_));
 sky130_fd_sc_hd__a2bb2oi_1 _16065_ (.A1_N(_06945_),
    .A2_N(net377),
    .B1(_05379_),
    .B2(_05393_),
    .Y(_05398_));
 sky130_fd_sc_hd__o22ai_4 _16066_ (.A1(_06945_),
    .A2(net377),
    .B1(_05378_),
    .B2(_05391_),
    .Y(_05399_));
 sky130_fd_sc_hd__o2bb2ai_2 _16067_ (.A1_N(_05176_),
    .A2_N(_05184_),
    .B1(_05394_),
    .B2(_07033_),
    .Y(_05400_));
 sky130_fd_sc_hd__o211ai_2 _16068_ (.A1(_05395_),
    .A2(_05378_),
    .B1(_05240_),
    .C1(_05399_),
    .Y(_05401_));
 sky130_fd_sc_hd__o21ai_2 _16069_ (.A1(_05396_),
    .A2(_05398_),
    .B1(_05238_),
    .Y(_05402_));
 sky130_fd_sc_hd__a2bb2oi_2 _16070_ (.A1_N(net328),
    .A2_N(_12681_),
    .B1(_05401_),
    .B2(_05402_),
    .Y(_05404_));
 sky130_fd_sc_hd__and3_1 _16071_ (.A(_12703_),
    .B(_05379_),
    .C(_05393_),
    .X(_05405_));
 sky130_fd_sc_hd__a21oi_4 _16072_ (.A1(_05379_),
    .A2(_05393_),
    .B1(net313),
    .Y(_05406_));
 sky130_fd_sc_hd__or3_1 _16073_ (.A(net328),
    .B(_12681_),
    .C(_05394_),
    .X(_05407_));
 sky130_fd_sc_hd__o221a_2 _16074_ (.A1(net328),
    .A2(_12681_),
    .B1(_05396_),
    .B2(_05400_),
    .C1(_05402_),
    .X(_05408_));
 sky130_fd_sc_hd__o221ai_4 _16075_ (.A1(net328),
    .A2(_12681_),
    .B1(_05396_),
    .B2(_05400_),
    .C1(_05402_),
    .Y(_05409_));
 sky130_fd_sc_hd__a31o_1 _16076_ (.A1(_05401_),
    .A2(_05402_),
    .A3(net313),
    .B1(_05406_),
    .X(_05410_));
 sky130_fd_sc_hd__or4_4 _16077_ (.A(net324),
    .B(net322),
    .C(_05404_),
    .D(_05405_),
    .X(_05411_));
 sky130_fd_sc_hd__a2bb2oi_4 _16078_ (.A1_N(net392),
    .A2_N(net382),
    .B1(_05407_),
    .B2(_05409_),
    .Y(_05412_));
 sky130_fd_sc_hd__o22ai_4 _16079_ (.A1(net392),
    .A2(net382),
    .B1(_05406_),
    .B2(_05408_),
    .Y(_05413_));
 sky130_fd_sc_hd__o221a_2 _16080_ (.A1(net380),
    .A2(net391),
    .B1(net313),
    .B2(_05394_),
    .C1(_05409_),
    .X(_05415_));
 sky130_fd_sc_hd__o221ai_4 _16081_ (.A1(net380),
    .A2(net391),
    .B1(net313),
    .B2(_05394_),
    .C1(_05409_),
    .Y(_05416_));
 sky130_fd_sc_hd__a22oi_4 _16082_ (.A1(_05173_),
    .A2(_05202_),
    .B1(_05204_),
    .B2(_05192_),
    .Y(_05417_));
 sky130_fd_sc_hd__o2bb2ai_4 _16083_ (.A1_N(_05173_),
    .A2_N(_05202_),
    .B1(_05193_),
    .B2(_05203_),
    .Y(_05418_));
 sky130_fd_sc_hd__o21ai_2 _16084_ (.A1(_05412_),
    .A2(_05415_),
    .B1(_05417_),
    .Y(_05419_));
 sky130_fd_sc_hd__nand3_2 _16085_ (.A(_05413_),
    .B(_05416_),
    .C(_05418_),
    .Y(_05420_));
 sky130_fd_sc_hd__o21ai_2 _16086_ (.A1(_05412_),
    .A2(_05415_),
    .B1(_05418_),
    .Y(_05421_));
 sky130_fd_sc_hd__nand2_1 _16087_ (.A(_05417_),
    .B(_05416_),
    .Y(_05422_));
 sky130_fd_sc_hd__o211ai_2 _16088_ (.A1(_06343_),
    .A2(_05410_),
    .B1(_05417_),
    .C1(_05413_),
    .Y(_05423_));
 sky130_fd_sc_hd__o221ai_2 _16089_ (.A1(net324),
    .A2(net322),
    .B1(_05412_),
    .B2(_05422_),
    .C1(_05421_),
    .Y(_05424_));
 sky130_fd_sc_hd__nand3_2 _16090_ (.A(_05419_),
    .B(_05420_),
    .C(net310),
    .Y(_05426_));
 sky130_fd_sc_hd__o221a_1 _16091_ (.A1(_14458_),
    .A2(_00000_),
    .B1(_05394_),
    .B2(net313),
    .C1(_05409_),
    .X(_05427_));
 sky130_fd_sc_hd__or4_1 _16092_ (.A(net324),
    .B(net322),
    .C(_05406_),
    .D(_05408_),
    .X(_05428_));
 sky130_fd_sc_hd__o31a_1 _16093_ (.A1(net310),
    .A2(_05406_),
    .A3(_05408_),
    .B1(_05426_),
    .X(_05429_));
 sky130_fd_sc_hd__nand4_2 _16094_ (.A(_03864_),
    .B(_03886_),
    .C(_05200_),
    .D(_05201_),
    .Y(_05430_));
 sky130_fd_sc_hd__a32oi_4 _16095_ (.A1(_05556_),
    .A2(_03864_),
    .A3(_03886_),
    .B1(_05208_),
    .B2(_05205_),
    .Y(_05431_));
 sky130_fd_sc_hd__o211ai_4 _16096_ (.A1(net386),
    .A2(_05206_),
    .B1(_05209_),
    .C1(_05430_),
    .Y(_05432_));
 sky130_fd_sc_hd__nand4_1 _16097_ (.A(_05209_),
    .B(_05214_),
    .C(_05430_),
    .D(_05851_),
    .Y(_05433_));
 sky130_fd_sc_hd__o21ai_1 _16098_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_05432_),
    .Y(_05434_));
 sky130_fd_sc_hd__a31o_1 _16099_ (.A1(_05434_),
    .A2(_01962_),
    .A3(_05433_),
    .B1(_05429_),
    .X(_05435_));
 sky130_fd_sc_hd__nand4_2 _16100_ (.A(_05429_),
    .B(_05433_),
    .C(_05434_),
    .D(_01962_),
    .Y(_05437_));
 sky130_fd_sc_hd__a311o_2 _16101_ (.A1(_05419_),
    .A2(_05420_),
    .A3(net310),
    .B1(_05427_),
    .C1(_01962_),
    .X(_05438_));
 sky130_fd_sc_hd__a311oi_1 _16102_ (.A1(_05419_),
    .A2(_05420_),
    .A3(net310),
    .B1(_05427_),
    .C1(_05851_),
    .Y(_05439_));
 sky130_fd_sc_hd__o211ai_2 _16103_ (.A1(net310),
    .A2(_05410_),
    .B1(_05426_),
    .C1(_05862_),
    .Y(_05440_));
 sky130_fd_sc_hd__a31oi_4 _16104_ (.A1(_05421_),
    .A2(_05423_),
    .A3(net310),
    .B1(_05862_),
    .Y(_05441_));
 sky130_fd_sc_hd__o211ai_1 _16105_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_05411_),
    .C1(_05424_),
    .Y(_05442_));
 sky130_fd_sc_hd__a32oi_4 _16106_ (.A1(_05862_),
    .A2(_05426_),
    .A3(_05428_),
    .B1(_05441_),
    .B2(_05411_),
    .Y(_05443_));
 sky130_fd_sc_hd__nand3_1 _16107_ (.A(_05432_),
    .B(_05440_),
    .C(_05442_),
    .Y(_05444_));
 sky130_fd_sc_hd__o221ai_4 _16108_ (.A1(net306),
    .A2(net303),
    .B1(_05432_),
    .B2(_05443_),
    .C1(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__nand2_2 _16109_ (.A(_05438_),
    .B(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__nand2_2 _16110_ (.A(_05435_),
    .B(_05437_),
    .Y(_05448_));
 sky130_fd_sc_hd__o32ai_4 _16111_ (.A1(_05250_),
    .A2(_05210_),
    .A3(_05212_),
    .B1(_03953_),
    .B2(_05219_),
    .Y(_05449_));
 sky130_fd_sc_hd__a21oi_2 _16112_ (.A1(_05217_),
    .A2(_05223_),
    .B1(net386),
    .Y(_05450_));
 sky130_fd_sc_hd__o21ai_4 _16113_ (.A1(net398),
    .A2(net397),
    .B1(_05449_),
    .Y(_05451_));
 sky130_fd_sc_hd__a221oi_4 _16114_ (.A1(_05512_),
    .A2(_05534_),
    .B1(_05220_),
    .B2(_03941_),
    .C1(_05216_),
    .Y(_05452_));
 sky130_fd_sc_hd__o221ai_4 _16115_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_03953_),
    .B2(_05219_),
    .C1(_05217_),
    .Y(_05453_));
 sky130_fd_sc_hd__o2111a_1 _16116_ (.A1(net301),
    .A2(net300),
    .B1(_05453_),
    .C1(_05446_),
    .D1(_05451_),
    .X(_05454_));
 sky130_fd_sc_hd__o2111ai_4 _16117_ (.A1(net301),
    .A2(net300),
    .B1(_05453_),
    .C1(_05446_),
    .D1(_05451_),
    .Y(_05455_));
 sky130_fd_sc_hd__a31oi_4 _16118_ (.A1(_05451_),
    .A2(_05453_),
    .A3(net275),
    .B1(_05446_),
    .Y(_05456_));
 sky130_fd_sc_hd__a31o_1 _16119_ (.A1(_05451_),
    .A2(_05453_),
    .A3(net275),
    .B1(_05446_),
    .X(_05457_));
 sky130_fd_sc_hd__nand3_1 _16120_ (.A(_05445_),
    .B(net386),
    .C(_05438_),
    .Y(_05459_));
 sky130_fd_sc_hd__nand3_1 _16121_ (.A(_05556_),
    .B(_05435_),
    .C(_05437_),
    .Y(_05460_));
 sky130_fd_sc_hd__o211ai_1 _16122_ (.A1(net386),
    .A2(_05448_),
    .B1(_05449_),
    .C1(_05459_),
    .Y(_05461_));
 sky130_fd_sc_hd__a21o_1 _16123_ (.A1(_05459_),
    .A2(_05460_),
    .B1(_05449_),
    .X(_05462_));
 sky130_fd_sc_hd__nand3_1 _16124_ (.A(_05462_),
    .B(net275),
    .C(_05461_),
    .Y(_05463_));
 sky130_fd_sc_hd__or3_1 _16125_ (.A(net301),
    .B(net300),
    .C(_05448_),
    .X(_05464_));
 sky130_fd_sc_hd__nor3_4 _16126_ (.A(_05250_),
    .B(_05454_),
    .C(_05456_),
    .Y(_05465_));
 sky130_fd_sc_hd__nand4_2 _16127_ (.A(_05207_),
    .B(_05229_),
    .C(_05455_),
    .D(_05457_),
    .Y(_05466_));
 sky130_fd_sc_hd__a21oi_2 _16128_ (.A1(_05455_),
    .A2(_05457_),
    .B1(net403),
    .Y(_05467_));
 sky130_fd_sc_hd__o21ai_1 _16129_ (.A1(_05454_),
    .A2(_05456_),
    .B1(_05250_),
    .Y(_05468_));
 sky130_fd_sc_hd__o21ai_1 _16130_ (.A1(_05465_),
    .A2(_05467_),
    .B1(_05225_),
    .Y(_05470_));
 sky130_fd_sc_hd__a31oi_4 _16131_ (.A1(_05250_),
    .A2(_05463_),
    .A3(_05464_),
    .B1(_05225_),
    .Y(_05471_));
 sky130_fd_sc_hd__nand4_1 _16132_ (.A(_05466_),
    .B(_05468_),
    .C(net1),
    .D(_05224_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand3_1 _16133_ (.A(_05470_),
    .B(_05472_),
    .C(net274),
    .Y(_05473_));
 sky130_fd_sc_hd__or4_1 _16134_ (.A(net297),
    .B(_05232_),
    .C(_05454_),
    .D(_05456_),
    .X(_05474_));
 sky130_fd_sc_hd__nand2_1 _16135_ (.A(_05473_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__inv_2 _16136_ (.A(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__or4_4 _16137_ (.A(net35),
    .B(net36),
    .C(net37),
    .D(_01908_),
    .X(_05477_));
 sky130_fd_sc_hd__o311a_4 _16138_ (.A1(net36),
    .A2(net37),
    .A3(_03975_),
    .B1(net38),
    .C1(net409),
    .X(_05478_));
 sky130_fd_sc_hd__a21oi_4 _16139_ (.A1(_05477_),
    .A2(net409),
    .B1(net38),
    .Y(_05479_));
 sky130_fd_sc_hd__and3b_4 _16140_ (.A_N(net38),
    .B(_05477_),
    .C(net409),
    .X(_05481_));
 sky130_fd_sc_hd__inv_2 _16141_ (.A(net270),
    .Y(_05482_));
 sky130_fd_sc_hd__a21boi_4 _16142_ (.A1(_05477_),
    .A2(net409),
    .B1_N(net38),
    .Y(_05483_));
 sky130_fd_sc_hd__inv_2 _16143_ (.A(net268),
    .Y(_05484_));
 sky130_fd_sc_hd__nor2_8 _16144_ (.A(_05478_),
    .B(_05479_),
    .Y(_05485_));
 sky130_fd_sc_hd__nor2_8 _16145_ (.A(net270),
    .B(net268),
    .Y(_05486_));
 sky130_fd_sc_hd__a21o_1 _16146_ (.A1(net1),
    .A2(_05485_),
    .B1(_05475_),
    .X(_05487_));
 sky130_fd_sc_hd__a21oi_1 _16147_ (.A1(_05473_),
    .A2(_05474_),
    .B1(_03289_),
    .Y(_05488_));
 sky130_fd_sc_hd__a21o_1 _16148_ (.A1(_05473_),
    .A2(_05474_),
    .B1(_03289_),
    .X(_05489_));
 sky130_fd_sc_hd__o31a_1 _16149_ (.A1(_03289_),
    .A2(_05476_),
    .A3(_05486_),
    .B1(_05487_),
    .X(_05490_));
 sky130_fd_sc_hd__inv_2 _16150_ (.A(_05490_),
    .Y(_05492_));
 sky130_fd_sc_hd__o21ai_1 _16151_ (.A1(_05051_),
    .A2(_05237_),
    .B1(_05490_),
    .Y(_05493_));
 sky130_fd_sc_hd__a311o_1 _16152_ (.A1(_02027_),
    .A2(_04063_),
    .A3(_05236_),
    .B1(_05490_),
    .C1(_05051_),
    .X(_05494_));
 sky130_fd_sc_hd__nand2_1 _16153_ (.A(_05493_),
    .B(_05494_),
    .Y(net70));
 sky130_fd_sc_hd__o2bb2a_1 _16154_ (.A1_N(_05237_),
    .A2_N(_05492_),
    .B1(_04832_),
    .B2(_04942_),
    .X(_05495_));
 sky130_fd_sc_hd__a21oi_4 _16155_ (.A1(_05417_),
    .A2(_05416_),
    .B1(_05412_),
    .Y(_05496_));
 sky130_fd_sc_hd__o32ai_4 _16156_ (.A1(_06332_),
    .A2(_05404_),
    .A3(_05405_),
    .B1(_05418_),
    .B2(_05415_),
    .Y(_05497_));
 sky130_fd_sc_hd__or4_4 _16157_ (.A(net4),
    .B(net5),
    .C(net6),
    .D(_02038_),
    .X(_05498_));
 sky130_fd_sc_hd__o21ai_4 _16158_ (.A1(net6),
    .A2(_05241_),
    .B1(net410),
    .Y(_05499_));
 sky130_fd_sc_hd__nor2_8 _16159_ (.A(net7),
    .B(_05499_),
    .Y(_05500_));
 sky130_fd_sc_hd__or3b_4 _16160_ (.A(_03399_),
    .B(net7),
    .C_N(_05498_),
    .X(_05502_));
 sky130_fd_sc_hd__and2_4 _16161_ (.A(_05499_),
    .B(net7),
    .X(_05503_));
 sky130_fd_sc_hd__nand2_8 _16162_ (.A(_05499_),
    .B(net7),
    .Y(_05504_));
 sky130_fd_sc_hd__o311a_4 _16163_ (.A1(net5),
    .A2(net6),
    .A3(_04150_),
    .B1(net7),
    .C1(net410),
    .X(_05505_));
 sky130_fd_sc_hd__a21oi_4 _16164_ (.A1(_05498_),
    .A2(net410),
    .B1(net7),
    .Y(_05506_));
 sky130_fd_sc_hd__nor2_8 _16165_ (.A(_05500_),
    .B(_05503_),
    .Y(_05507_));
 sky130_fd_sc_hd__nor2_2 _16166_ (.A(_05505_),
    .B(_05506_),
    .Y(_05508_));
 sky130_fd_sc_hd__or3_2 _16167_ (.A(_03178_),
    .B(_05505_),
    .C(_05506_),
    .X(_05509_));
 sky130_fd_sc_hd__o221a_1 _16168_ (.A1(net408),
    .A2(_05152_),
    .B1(_05500_),
    .B2(_05503_),
    .C1(net33),
    .X(_05510_));
 sky130_fd_sc_hd__a211o_1 _16169_ (.A1(net291),
    .A2(net33),
    .B1(_05242_),
    .C1(net317),
    .X(_05511_));
 sky130_fd_sc_hd__o31a_1 _16170_ (.A1(_05252_),
    .A2(_05505_),
    .A3(_05506_),
    .B1(_05511_),
    .X(_05513_));
 sky130_fd_sc_hd__o21ai_2 _16171_ (.A1(_05252_),
    .A2(net267),
    .B1(_05511_),
    .Y(_05514_));
 sky130_fd_sc_hd__o22ai_4 _16172_ (.A1(_04249_),
    .A2(net295),
    .B1(_05257_),
    .B2(_05254_),
    .Y(_05515_));
 sky130_fd_sc_hd__a21oi_1 _16173_ (.A1(_05256_),
    .A2(_05258_),
    .B1(_05514_),
    .Y(_05516_));
 sky130_fd_sc_hd__nand2_2 _16174_ (.A(_05515_),
    .B(_05513_),
    .Y(_05517_));
 sky130_fd_sc_hd__o221ai_4 _16175_ (.A1(_04249_),
    .A2(net295),
    .B1(_05257_),
    .B2(_05254_),
    .C1(_05514_),
    .Y(_05518_));
 sky130_fd_sc_hd__o21ai_1 _16176_ (.A1(_05513_),
    .A2(_05515_),
    .B1(_05174_),
    .Y(_05519_));
 sky130_fd_sc_hd__nand2_1 _16177_ (.A(_05517_),
    .B(_05518_),
    .Y(_05520_));
 sky130_fd_sc_hd__o32a_1 _16178_ (.A1(_03178_),
    .A2(_05505_),
    .A3(_05506_),
    .B1(net408),
    .B2(_05152_),
    .X(_05521_));
 sky130_fd_sc_hd__a22o_1 _16179_ (.A1(_05141_),
    .A2(_05163_),
    .B1(net291),
    .B2(net33),
    .X(_05522_));
 sky130_fd_sc_hd__o32a_4 _16180_ (.A1(_03178_),
    .A2(_05174_),
    .A3(net267),
    .B1(_05516_),
    .B2(_05519_),
    .X(_05524_));
 sky130_fd_sc_hd__o22ai_1 _16181_ (.A1(_05174_),
    .A2(_05509_),
    .B1(_05516_),
    .B2(_05519_),
    .Y(_05525_));
 sky130_fd_sc_hd__or3_4 _16182_ (.A(net402),
    .B(net400),
    .C(_05524_),
    .X(_05526_));
 sky130_fd_sc_hd__a311oi_4 _16183_ (.A1(_05517_),
    .A2(_05518_),
    .A3(_05174_),
    .B1(net298),
    .C1(_05510_),
    .Y(_05527_));
 sky130_fd_sc_hd__a311o_1 _16184_ (.A1(_05517_),
    .A2(_05518_),
    .A3(_05174_),
    .B1(net298),
    .C1(_05510_),
    .X(_05528_));
 sky130_fd_sc_hd__a22oi_4 _16185_ (.A1(_04173_),
    .A2(_04195_),
    .B1(_05520_),
    .B2(_05174_),
    .Y(_05529_));
 sky130_fd_sc_hd__a31o_1 _16186_ (.A1(_05141_),
    .A2(_05163_),
    .A3(_05520_),
    .B1(net299),
    .X(_05530_));
 sky130_fd_sc_hd__o21ai_2 _16187_ (.A1(net339),
    .A2(_04184_),
    .B1(_05525_),
    .Y(_05531_));
 sky130_fd_sc_hd__a21oi_4 _16188_ (.A1(_05529_),
    .A2(_05522_),
    .B1(_05527_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand2_1 _16189_ (.A(_05528_),
    .B(_05531_),
    .Y(_05533_));
 sky130_fd_sc_hd__a31oi_1 _16190_ (.A1(_05274_),
    .A2(_04569_),
    .A3(_04536_),
    .B1(_05269_),
    .Y(_05535_));
 sky130_fd_sc_hd__o2bb2ai_2 _16191_ (.A1_N(_02137_),
    .A2_N(_05264_),
    .B1(_05275_),
    .B2(_04591_),
    .Y(_05536_));
 sky130_fd_sc_hd__a21oi_1 _16192_ (.A1(_05277_),
    .A2(_04625_),
    .B1(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__o21bai_4 _16193_ (.A1(_05536_),
    .A2(_05279_),
    .B1_N(_05267_),
    .Y(_05538_));
 sky130_fd_sc_hd__a21oi_2 _16194_ (.A1(_05535_),
    .A2(_05280_),
    .B1(_05267_),
    .Y(_05539_));
 sky130_fd_sc_hd__a21oi_2 _16195_ (.A1(_05268_),
    .A2(_05284_),
    .B1(_05533_),
    .Y(_05540_));
 sky130_fd_sc_hd__o21ai_4 _16196_ (.A1(_05267_),
    .A2(_05537_),
    .B1(_05532_),
    .Y(_05541_));
 sky130_fd_sc_hd__o22ai_4 _16197_ (.A1(net402),
    .A2(net400),
    .B1(_05532_),
    .B2(_05538_),
    .Y(_05542_));
 sky130_fd_sc_hd__o221ai_4 _16198_ (.A1(net402),
    .A2(net400),
    .B1(_05532_),
    .B2(_05538_),
    .C1(_05541_),
    .Y(_05543_));
 sky130_fd_sc_hd__o22a_1 _16199_ (.A1(net388),
    .A2(_05524_),
    .B1(_05540_),
    .B2(_05542_),
    .X(_05544_));
 sky130_fd_sc_hd__o22ai_4 _16200_ (.A1(net388),
    .A2(_05524_),
    .B1(_05540_),
    .B2(_05542_),
    .Y(_05546_));
 sky130_fd_sc_hd__o2bb2ai_1 _16201_ (.A1_N(net319),
    .A2_N(_05288_),
    .B1(_05291_),
    .B2(_04734_),
    .Y(_05547_));
 sky130_fd_sc_hd__a22oi_2 _16202_ (.A1(_05265_),
    .A2(_05295_),
    .B1(_05299_),
    .B2(_05293_),
    .Y(_05548_));
 sky130_fd_sc_hd__o21ai_2 _16203_ (.A1(_05292_),
    .A2(_05298_),
    .B1(_05297_),
    .Y(_05549_));
 sky130_fd_sc_hd__a2bb2oi_4 _16204_ (.A1_N(_02049_),
    .A2_N(net342),
    .B1(_05526_),
    .B2(_05543_),
    .Y(_05550_));
 sky130_fd_sc_hd__o21ai_1 _16205_ (.A1(_02049_),
    .A2(net342),
    .B1(_05546_),
    .Y(_05551_));
 sky130_fd_sc_hd__o221a_1 _16206_ (.A1(net388),
    .A2(_05524_),
    .B1(_05540_),
    .B2(_05542_),
    .C1(_02137_),
    .X(_05552_));
 sky130_fd_sc_hd__nand3_4 _16207_ (.A(_05543_),
    .B(_02137_),
    .C(_05526_),
    .Y(_05553_));
 sky130_fd_sc_hd__nand3_1 _16208_ (.A(_05549_),
    .B(_05551_),
    .C(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__o21ai_1 _16209_ (.A1(_05550_),
    .A2(_05552_),
    .B1(_05548_),
    .Y(_05555_));
 sky130_fd_sc_hd__nand3_1 _16210_ (.A(_05555_),
    .B(net359),
    .C(_05554_),
    .Y(_05557_));
 sky130_fd_sc_hd__a211o_1 _16211_ (.A1(_05526_),
    .A2(_05543_),
    .B1(net384),
    .C1(net383),
    .X(_05558_));
 sky130_fd_sc_hd__o211ai_4 _16212_ (.A1(_05292_),
    .A2(_05298_),
    .B1(_05553_),
    .C1(_05297_),
    .Y(_05559_));
 sky130_fd_sc_hd__o2bb2ai_1 _16213_ (.A1_N(_05297_),
    .A2_N(_05547_),
    .B1(_05550_),
    .B2(_05552_),
    .Y(_05560_));
 sky130_fd_sc_hd__o211ai_4 _16214_ (.A1(_05550_),
    .A2(_05559_),
    .B1(net359),
    .C1(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__o21ai_2 _16215_ (.A1(net359),
    .A2(_05544_),
    .B1(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__and3_1 _16216_ (.A(_05562_),
    .B(_06826_),
    .C(_06804_),
    .X(_05563_));
 sky130_fd_sc_hd__a211o_2 _16217_ (.A1(_05558_),
    .A2(_05561_),
    .B1(net379),
    .C1(net378),
    .X(_05564_));
 sky130_fd_sc_hd__a2bb2oi_1 _16218_ (.A1_N(_00174_),
    .A2_N(_00196_),
    .B1(_05558_),
    .B2(_05561_),
    .Y(_05565_));
 sky130_fd_sc_hd__o211ai_4 _16219_ (.A1(_05546_),
    .A2(net359),
    .B1(net319),
    .C1(_05557_),
    .Y(_05566_));
 sky130_fd_sc_hd__o211a_1 _16220_ (.A1(net359),
    .A2(_05544_),
    .B1(net320),
    .C1(_05561_),
    .X(_05568_));
 sky130_fd_sc_hd__nand3_4 _16221_ (.A(_05561_),
    .B(net320),
    .C(_05558_),
    .Y(_05569_));
 sky130_fd_sc_hd__nand2_4 _16222_ (.A(_05566_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__o21ai_2 _16223_ (.A1(_04866_),
    .A2(_05309_),
    .B1(_05315_),
    .Y(_05571_));
 sky130_fd_sc_hd__a21oi_4 _16224_ (.A1(_05311_),
    .A2(_05313_),
    .B1(_05314_),
    .Y(_05572_));
 sky130_fd_sc_hd__a22oi_2 _16225_ (.A1(_05566_),
    .A2(_05569_),
    .B1(_05571_),
    .B2(_05313_),
    .Y(_05573_));
 sky130_fd_sc_hd__nand2_2 _16226_ (.A(_05570_),
    .B(_05572_),
    .Y(_05574_));
 sky130_fd_sc_hd__o2111a_1 _16227_ (.A1(net325),
    .A2(_05307_),
    .B1(_05566_),
    .C1(_05569_),
    .D1(_05571_),
    .X(_05575_));
 sky130_fd_sc_hd__o2111ai_4 _16228_ (.A1(net325),
    .A2(_05307_),
    .B1(_05566_),
    .C1(_05569_),
    .D1(_05571_),
    .Y(_05576_));
 sky130_fd_sc_hd__o211ai_4 _16229_ (.A1(_05570_),
    .A2(_05572_),
    .B1(net357),
    .C1(_05574_),
    .Y(_05577_));
 sky130_fd_sc_hd__o22ai_2 _16230_ (.A1(net379),
    .A2(net378),
    .B1(_05573_),
    .B2(_05575_),
    .Y(_05579_));
 sky130_fd_sc_hd__o31a_1 _16231_ (.A1(_06848_),
    .A2(_05573_),
    .A3(_05575_),
    .B1(_05564_),
    .X(_05580_));
 sky130_fd_sc_hd__a311o_1 _16232_ (.A1(_05574_),
    .A2(_05576_),
    .A3(net357),
    .B1(net356),
    .C1(_05563_),
    .X(_05581_));
 sky130_fd_sc_hd__a21oi_2 _16233_ (.A1(_05324_),
    .A2(net330),
    .B1(_05332_),
    .Y(_05582_));
 sky130_fd_sc_hd__o21ai_4 _16234_ (.A1(_05040_),
    .A2(_05331_),
    .B1(_05328_),
    .Y(_05583_));
 sky130_fd_sc_hd__a21oi_1 _16235_ (.A1(_05325_),
    .A2(net331),
    .B1(_05333_),
    .Y(_05584_));
 sky130_fd_sc_hd__a311oi_4 _16236_ (.A1(_05574_),
    .A2(_05576_),
    .A3(net357),
    .B1(net325),
    .C1(_05563_),
    .Y(_05585_));
 sky130_fd_sc_hd__o211ai_4 _16237_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_05564_),
    .C1(_05577_),
    .Y(_05586_));
 sky130_fd_sc_hd__a2bb2oi_4 _16238_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_05564_),
    .B2(_05577_),
    .Y(_05587_));
 sky130_fd_sc_hd__o211ai_2 _16239_ (.A1(net357),
    .A2(_05562_),
    .B1(_05579_),
    .C1(net325),
    .Y(_05588_));
 sky130_fd_sc_hd__o211ai_1 _16240_ (.A1(_05329_),
    .A2(_05582_),
    .B1(_05586_),
    .C1(_05588_),
    .Y(_05590_));
 sky130_fd_sc_hd__o22ai_1 _16241_ (.A1(_05327_),
    .A2(_05584_),
    .B1(_05585_),
    .B2(_05587_),
    .Y(_05591_));
 sky130_fd_sc_hd__nand3_1 _16242_ (.A(_05590_),
    .B(_05591_),
    .C(net356),
    .Y(_05592_));
 sky130_fd_sc_hd__o311a_2 _16243_ (.A1(net379),
    .A2(net378),
    .A3(_05562_),
    .B1(_05579_),
    .C1(_07724_),
    .X(_05593_));
 sky130_fd_sc_hd__o2111ai_4 _16244_ (.A1(net330),
    .A2(_05324_),
    .B1(_05583_),
    .C1(_05586_),
    .D1(_05588_),
    .Y(_05594_));
 sky130_fd_sc_hd__o22ai_4 _16245_ (.A1(_05329_),
    .A2(_05582_),
    .B1(_05585_),
    .B2(_05587_),
    .Y(_05595_));
 sky130_fd_sc_hd__o211ai_2 _16246_ (.A1(net372),
    .A2(net371),
    .B1(_05594_),
    .C1(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__a31o_2 _16247_ (.A1(_05594_),
    .A2(_05595_),
    .A3(net356),
    .B1(_05593_),
    .X(_05597_));
 sky130_fd_sc_hd__a31oi_4 _16248_ (.A1(_05594_),
    .A2(_05595_),
    .A3(net356),
    .B1(_05593_),
    .Y(_05598_));
 sky130_fd_sc_hd__and3_1 _16249_ (.A(_05597_),
    .B(_11287_),
    .C(_11265_),
    .X(_05599_));
 sky130_fd_sc_hd__o211ai_4 _16250_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_05581_),
    .C1(_05592_),
    .Y(_05601_));
 sky130_fd_sc_hd__a31o_1 _16251_ (.A1(_05594_),
    .A2(_05595_),
    .A3(net356),
    .B1(net330),
    .X(_05602_));
 sky130_fd_sc_hd__o211a_1 _16252_ (.A1(net356),
    .A2(_05580_),
    .B1(net331),
    .C1(_05596_),
    .X(_05603_));
 sky130_fd_sc_hd__o211ai_4 _16253_ (.A1(net356),
    .A2(_05580_),
    .B1(net331),
    .C1(_05596_),
    .Y(_05604_));
 sky130_fd_sc_hd__a21oi_1 _16254_ (.A1(net348),
    .A2(_05342_),
    .B1(_05351_),
    .Y(_05605_));
 sky130_fd_sc_hd__o21ai_1 _16255_ (.A1(_05349_),
    .A2(_05350_),
    .B1(_05346_),
    .Y(_05606_));
 sky130_fd_sc_hd__o22ai_4 _16256_ (.A1(_05334_),
    .A2(_05347_),
    .B1(_05351_),
    .B2(_05345_),
    .Y(_05607_));
 sky130_fd_sc_hd__o2111ai_1 _16257_ (.A1(_05349_),
    .A2(_05350_),
    .B1(_05601_),
    .C1(_05604_),
    .D1(_05346_),
    .Y(_05608_));
 sky130_fd_sc_hd__a21o_1 _16258_ (.A1(_05601_),
    .A2(_05604_),
    .B1(_05607_),
    .X(_05609_));
 sky130_fd_sc_hd__nand3_2 _16259_ (.A(_05609_),
    .B(_08721_),
    .C(_05608_),
    .Y(_05610_));
 sky130_fd_sc_hd__or3_1 _16260_ (.A(net353),
    .B(net352),
    .C(_05598_),
    .X(_05612_));
 sky130_fd_sc_hd__o2bb2ai_1 _16261_ (.A1_N(_05601_),
    .A2_N(_05604_),
    .B1(_05605_),
    .B2(_05349_),
    .Y(_05613_));
 sky130_fd_sc_hd__nand3_1 _16262_ (.A(_05606_),
    .B(_05604_),
    .C(_05601_),
    .Y(_05614_));
 sky130_fd_sc_hd__nand3_2 _16263_ (.A(_05613_),
    .B(_05614_),
    .C(_08721_),
    .Y(_05615_));
 sky130_fd_sc_hd__o21ai_2 _16264_ (.A1(_08721_),
    .A2(_05597_),
    .B1(_05610_),
    .Y(_05616_));
 sky130_fd_sc_hd__o21ai_1 _16265_ (.A1(_09763_),
    .A2(_09774_),
    .B1(_05616_),
    .Y(_05617_));
 sky130_fd_sc_hd__a2bb2oi_2 _16266_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_05612_),
    .B2(_05615_),
    .Y(_05618_));
 sky130_fd_sc_hd__o211ai_4 _16267_ (.A1(_08721_),
    .A2(_05597_),
    .B1(_05610_),
    .C1(net348),
    .Y(_05619_));
 sky130_fd_sc_hd__o221a_4 _16268_ (.A1(_09971_),
    .A2(net363),
    .B1(_05598_),
    .B2(_08721_),
    .C1(_05615_),
    .X(_05620_));
 sky130_fd_sc_hd__o221ai_4 _16269_ (.A1(_09971_),
    .A2(net363),
    .B1(_05598_),
    .B2(_08721_),
    .C1(_05615_),
    .Y(_05621_));
 sky130_fd_sc_hd__a32oi_4 _16270_ (.A1(_05360_),
    .A2(_08907_),
    .A3(_05356_),
    .B1(_05142_),
    .B2(_05151_),
    .Y(_05622_));
 sky130_fd_sc_hd__o2bb2ai_1 _16271_ (.A1_N(_05142_),
    .A2_N(_05151_),
    .B1(_08918_),
    .B2(_05361_),
    .Y(_05623_));
 sky130_fd_sc_hd__o21ai_1 _16272_ (.A1(_08907_),
    .A2(_05362_),
    .B1(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__a21oi_2 _16273_ (.A1(_05364_),
    .A2(_05371_),
    .B1(_05372_),
    .Y(_05625_));
 sky130_fd_sc_hd__o211ai_4 _16274_ (.A1(_05372_),
    .A2(_05622_),
    .B1(_05621_),
    .C1(_05619_),
    .Y(_05626_));
 sky130_fd_sc_hd__o21ai_4 _16275_ (.A1(_05618_),
    .A2(_05620_),
    .B1(_05625_),
    .Y(_05627_));
 sky130_fd_sc_hd__o21ai_1 _16276_ (.A1(_05618_),
    .A2(_05620_),
    .B1(_05624_),
    .Y(_05628_));
 sky130_fd_sc_hd__o2111ai_1 _16277_ (.A1(_05362_),
    .A2(_08907_),
    .B1(_05621_),
    .C1(_05619_),
    .D1(_05623_),
    .Y(_05629_));
 sky130_fd_sc_hd__nand3_1 _16278_ (.A(_05628_),
    .B(_05629_),
    .C(net337),
    .Y(_05630_));
 sky130_fd_sc_hd__o211a_1 _16279_ (.A1(_08721_),
    .A2(_05597_),
    .B1(_05610_),
    .C1(_09840_),
    .X(_05631_));
 sky130_fd_sc_hd__or3_1 _16280_ (.A(net350),
    .B(net349),
    .C(_05616_),
    .X(_05633_));
 sky130_fd_sc_hd__o211ai_4 _16281_ (.A1(net350),
    .A2(net349),
    .B1(_05626_),
    .C1(_05627_),
    .Y(_05634_));
 sky130_fd_sc_hd__and3_2 _16282_ (.A(_11079_),
    .B(_05617_),
    .C(_05630_),
    .X(_05635_));
 sky130_fd_sc_hd__a211o_2 _16283_ (.A1(_05633_),
    .A2(_05634_),
    .B1(net347),
    .C1(net346),
    .X(_05636_));
 sky130_fd_sc_hd__o211a_1 _16284_ (.A1(_04117_),
    .A2(_05160_),
    .B1(_05164_),
    .C1(_05388_),
    .X(_05637_));
 sky130_fd_sc_hd__a22oi_4 _16285_ (.A1(_05384_),
    .A2(_05377_),
    .B1(_05383_),
    .B2(_05388_),
    .Y(_05638_));
 sky130_fd_sc_hd__a311oi_4 _16286_ (.A1(_05627_),
    .A2(net337),
    .A3(_05626_),
    .B1(_05631_),
    .C1(_08918_),
    .Y(_05639_));
 sky130_fd_sc_hd__o211ai_4 _16287_ (.A1(net337),
    .A2(_05616_),
    .B1(_08907_),
    .C1(_05634_),
    .Y(_05640_));
 sky130_fd_sc_hd__a2bb2oi_2 _16288_ (.A1_N(_08819_),
    .A2_N(net367),
    .B1(_05633_),
    .B2(_05634_),
    .Y(_05641_));
 sky130_fd_sc_hd__o211ai_2 _16289_ (.A1(_08819_),
    .A2(net367),
    .B1(_05617_),
    .C1(_05630_),
    .Y(_05642_));
 sky130_fd_sc_hd__nand3_4 _16290_ (.A(_05638_),
    .B(_05640_),
    .C(_05642_),
    .Y(_05644_));
 sky130_fd_sc_hd__o22ai_4 _16291_ (.A1(_05385_),
    .A2(_05637_),
    .B1(_05639_),
    .B2(_05641_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand3_4 _16292_ (.A(_05645_),
    .B(net334),
    .C(_05644_),
    .Y(_05646_));
 sky130_fd_sc_hd__a31oi_4 _16293_ (.A1(_05645_),
    .A2(net334),
    .A3(_05644_),
    .B1(_05635_),
    .Y(_05647_));
 sky130_fd_sc_hd__a21oi_4 _16294_ (.A1(_05636_),
    .A2(_05646_),
    .B1(net313),
    .Y(_05648_));
 sky130_fd_sc_hd__or3_2 _16295_ (.A(net328),
    .B(_12681_),
    .C(_05647_),
    .X(_05649_));
 sky130_fd_sc_hd__o21ai_4 _16296_ (.A1(_07033_),
    .A2(_05394_),
    .B1(_05238_),
    .Y(_05650_));
 sky130_fd_sc_hd__o21ai_1 _16297_ (.A1(_05238_),
    .A2(_05396_),
    .B1(_05399_),
    .Y(_05651_));
 sky130_fd_sc_hd__a311oi_4 _16298_ (.A1(_05645_),
    .A2(net334),
    .A3(_05644_),
    .B1(_05635_),
    .C1(_07899_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand3_4 _16299_ (.A(_05646_),
    .B(_07888_),
    .C(_05636_),
    .Y(_05653_));
 sky130_fd_sc_hd__a2bb2oi_2 _16300_ (.A1_N(net389),
    .A2_N(net370),
    .B1(_05636_),
    .B2(_05646_),
    .Y(_05655_));
 sky130_fd_sc_hd__a22o_2 _16301_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_05636_),
    .B2(_05646_),
    .X(_05656_));
 sky130_fd_sc_hd__o211ai_4 _16302_ (.A1(_05395_),
    .A2(_05378_),
    .B1(_05653_),
    .C1(_05650_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand3_4 _16303_ (.A(_05656_),
    .B(_05651_),
    .C(_05653_),
    .Y(_05658_));
 sky130_fd_sc_hd__o2bb2ai_4 _16304_ (.A1_N(_05397_),
    .A2_N(_05650_),
    .B1(_05652_),
    .B2(_05655_),
    .Y(_05659_));
 sky130_fd_sc_hd__o211a_1 _16305_ (.A1(_05655_),
    .A2(_05657_),
    .B1(net313),
    .C1(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__o211ai_2 _16306_ (.A1(_05655_),
    .A2(_05657_),
    .B1(net313),
    .C1(_05659_),
    .Y(_05661_));
 sky130_fd_sc_hd__a31oi_4 _16307_ (.A1(_05658_),
    .A2(_05659_),
    .A3(net313),
    .B1(_05648_),
    .Y(_05662_));
 sky130_fd_sc_hd__a31o_4 _16308_ (.A1(_05658_),
    .A2(_05659_),
    .A3(net313),
    .B1(_05648_),
    .X(_05663_));
 sky130_fd_sc_hd__a31oi_1 _16309_ (.A1(_05658_),
    .A2(_05659_),
    .A3(net313),
    .B1(_07044_),
    .Y(_05664_));
 sky130_fd_sc_hd__o21ai_1 _16310_ (.A1(_06989_),
    .A2(_07011_),
    .B1(_05661_),
    .Y(_05666_));
 sky130_fd_sc_hd__a311oi_4 _16311_ (.A1(_05658_),
    .A2(_05659_),
    .A3(net313),
    .B1(_05648_),
    .C1(_07044_),
    .Y(_05667_));
 sky130_fd_sc_hd__a22oi_4 _16312_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_05649_),
    .B2(_05661_),
    .Y(_05668_));
 sky130_fd_sc_hd__o22ai_4 _16313_ (.A1(_06945_),
    .A2(net377),
    .B1(_05648_),
    .B2(_05660_),
    .Y(_05669_));
 sky130_fd_sc_hd__a221oi_2 _16314_ (.A1(_05664_),
    .A2(_05649_),
    .B1(_05422_),
    .B2(_05413_),
    .C1(_05668_),
    .Y(_05670_));
 sky130_fd_sc_hd__o211ai_4 _16315_ (.A1(_05666_),
    .A2(_05648_),
    .B1(_05497_),
    .C1(_05669_),
    .Y(_05671_));
 sky130_fd_sc_hd__o21a_1 _16316_ (.A1(_05667_),
    .A2(_05668_),
    .B1(_05496_),
    .X(_05672_));
 sky130_fd_sc_hd__o21ai_4 _16317_ (.A1(_05667_),
    .A2(_05668_),
    .B1(_05496_),
    .Y(_05673_));
 sky130_fd_sc_hd__o22ai_4 _16318_ (.A1(net324),
    .A2(net322),
    .B1(_05670_),
    .B2(_05672_),
    .Y(_05674_));
 sky130_fd_sc_hd__and3_1 _16319_ (.A(_00022_),
    .B(_00044_),
    .C(_05663_),
    .X(_05675_));
 sky130_fd_sc_hd__or3_1 _16320_ (.A(net324),
    .B(net322),
    .C(_05662_),
    .X(_05677_));
 sky130_fd_sc_hd__nand3_4 _16321_ (.A(_05673_),
    .B(net310),
    .C(_05671_),
    .Y(_05678_));
 sky130_fd_sc_hd__a31o_1 _16322_ (.A1(_05673_),
    .A2(net310),
    .A3(_05671_),
    .B1(_05675_),
    .X(_05679_));
 sky130_fd_sc_hd__o31a_1 _16323_ (.A1(net324),
    .A2(net322),
    .A3(_05662_),
    .B1(_05678_),
    .X(_05680_));
 sky130_fd_sc_hd__o311a_1 _16324_ (.A1(net324),
    .A2(_05663_),
    .A3(net322),
    .B1(_01973_),
    .C1(_05674_),
    .X(_05681_));
 sky130_fd_sc_hd__or3_2 _16325_ (.A(net305),
    .B(net303),
    .C(_05680_),
    .X(_05682_));
 sky130_fd_sc_hd__a2bb2oi_2 _16326_ (.A1_N(net393),
    .A2_N(net382),
    .B1(_05677_),
    .B2(_05678_),
    .Y(_05683_));
 sky130_fd_sc_hd__o211ai_4 _16327_ (.A1(_05663_),
    .A2(net310),
    .B1(_06343_),
    .C1(_05674_),
    .Y(_05684_));
 sky130_fd_sc_hd__o221a_1 _16328_ (.A1(_06289_),
    .A2(net391),
    .B1(net310),
    .B2(_05662_),
    .C1(_05678_),
    .X(_05685_));
 sky130_fd_sc_hd__o221ai_4 _16329_ (.A1(_06289_),
    .A2(net391),
    .B1(net310),
    .B2(_05662_),
    .C1(_05678_),
    .Y(_05686_));
 sky130_fd_sc_hd__o21ai_1 _16330_ (.A1(_05432_),
    .A2(_05439_),
    .B1(_05442_),
    .Y(_05688_));
 sky130_fd_sc_hd__a22oi_4 _16331_ (.A1(_05411_),
    .A2(_05441_),
    .B1(_05440_),
    .B2(_05431_),
    .Y(_05689_));
 sky130_fd_sc_hd__nand3_2 _16332_ (.A(_05684_),
    .B(_05686_),
    .C(_05688_),
    .Y(_05690_));
 sky130_fd_sc_hd__o21ai_2 _16333_ (.A1(_05683_),
    .A2(_05685_),
    .B1(_05689_),
    .Y(_05691_));
 sky130_fd_sc_hd__o21bai_2 _16334_ (.A1(_05683_),
    .A2(_05685_),
    .B1_N(_05689_),
    .Y(_05692_));
 sky130_fd_sc_hd__o21ai_2 _16335_ (.A1(_06343_),
    .A2(_05679_),
    .B1(_05689_),
    .Y(_05693_));
 sky130_fd_sc_hd__nand3_2 _16336_ (.A(_05684_),
    .B(_05686_),
    .C(_05689_),
    .Y(_05694_));
 sky130_fd_sc_hd__nand3_2 _16337_ (.A(_05691_),
    .B(_01962_),
    .C(_05690_),
    .Y(_05695_));
 sky130_fd_sc_hd__o221a_1 _16338_ (.A1(_01919_),
    .A2(_01930_),
    .B1(_05662_),
    .B2(net310),
    .C1(_05678_),
    .X(_05696_));
 sky130_fd_sc_hd__a311o_2 _16339_ (.A1(_05673_),
    .A2(net310),
    .A3(_05671_),
    .B1(_05675_),
    .C1(_01962_),
    .X(_05697_));
 sky130_fd_sc_hd__a31o_1 _16340_ (.A1(_05691_),
    .A2(_01962_),
    .A3(_05690_),
    .B1(_05696_),
    .X(_05699_));
 sky130_fd_sc_hd__a31o_1 _16341_ (.A1(_05692_),
    .A2(_05694_),
    .A3(_01962_),
    .B1(_05681_),
    .X(_05700_));
 sky130_fd_sc_hd__a32oi_4 _16342_ (.A1(_05223_),
    .A2(net386),
    .A3(_05217_),
    .B1(_05438_),
    .B2(_05445_),
    .Y(_05701_));
 sky130_fd_sc_hd__a21oi_1 _16343_ (.A1(_05446_),
    .A2(_05453_),
    .B1(_05450_),
    .Y(_05702_));
 sky130_fd_sc_hd__o21ai_2 _16344_ (.A1(_05448_),
    .A2(_05452_),
    .B1(_05451_),
    .Y(_05703_));
 sky130_fd_sc_hd__o211a_1 _16345_ (.A1(_05448_),
    .A2(_05452_),
    .B1(_05451_),
    .C1(_05851_),
    .X(_05704_));
 sky130_fd_sc_hd__o211ai_2 _16346_ (.A1(_05448_),
    .A2(_05452_),
    .B1(_05451_),
    .C1(_05851_),
    .Y(_05705_));
 sky130_fd_sc_hd__o22a_1 _16347_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_05450_),
    .B2(_05701_),
    .X(_05706_));
 sky130_fd_sc_hd__o22ai_2 _16348_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_05450_),
    .B2(_05701_),
    .Y(_05707_));
 sky130_fd_sc_hd__a31o_2 _16349_ (.A1(_05707_),
    .A2(net275),
    .A3(_05705_),
    .B1(_05700_),
    .X(_05708_));
 sky130_fd_sc_hd__nand4_4 _16350_ (.A(_05700_),
    .B(_05705_),
    .C(_05707_),
    .D(net275),
    .Y(_05710_));
 sky130_fd_sc_hd__a31oi_4 _16351_ (.A1(_05692_),
    .A2(_05694_),
    .A3(_01962_),
    .B1(_05862_),
    .Y(_05711_));
 sky130_fd_sc_hd__a311o_1 _16352_ (.A1(_05692_),
    .A2(_05694_),
    .A3(_01962_),
    .B1(_05681_),
    .C1(_05862_),
    .X(_05712_));
 sky130_fd_sc_hd__a311oi_1 _16353_ (.A1(_05691_),
    .A2(_01962_),
    .A3(_05690_),
    .B1(_05696_),
    .C1(_05851_),
    .Y(_05713_));
 sky130_fd_sc_hd__o211ai_2 _16354_ (.A1(_01962_),
    .A2(_05679_),
    .B1(_05695_),
    .C1(_05862_),
    .Y(_05714_));
 sky130_fd_sc_hd__o211ai_2 _16355_ (.A1(_05450_),
    .A2(_05701_),
    .B1(_05712_),
    .C1(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__a32oi_4 _16356_ (.A1(_05862_),
    .A2(_05695_),
    .A3(_05697_),
    .B1(_05711_),
    .B2(_05682_),
    .Y(_05716_));
 sky130_fd_sc_hd__o221ai_4 _16357_ (.A1(net301),
    .A2(net300),
    .B1(_05703_),
    .B2(_05716_),
    .C1(_05715_),
    .Y(_05717_));
 sky130_fd_sc_hd__o41a_1 _16358_ (.A1(_04040_),
    .A2(_05699_),
    .A3(_05704_),
    .A4(_05706_),
    .B1(_05708_),
    .X(_05718_));
 sky130_fd_sc_hd__nand2_4 _16359_ (.A(_05708_),
    .B(_05710_),
    .Y(_05719_));
 sky130_fd_sc_hd__a31oi_1 _16360_ (.A1(_05468_),
    .A2(_05224_),
    .A3(net1),
    .B1(_05465_),
    .Y(_05721_));
 sky130_fd_sc_hd__o21ai_1 _16361_ (.A1(_05225_),
    .A2(_05467_),
    .B1(_05466_),
    .Y(_05722_));
 sky130_fd_sc_hd__o221ai_4 _16362_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_05225_),
    .B2(_05467_),
    .C1(_05466_),
    .Y(_05723_));
 sky130_fd_sc_hd__o22ai_2 _16363_ (.A1(net398),
    .A2(net397),
    .B1(_05465_),
    .B2(_05471_),
    .Y(_05724_));
 sky130_fd_sc_hd__o2111ai_4 _16364_ (.A1(net297),
    .A2(_05232_),
    .B1(_05718_),
    .C1(_05723_),
    .D1(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__a31o_1 _16365_ (.A1(_05724_),
    .A2(net274),
    .A3(_05723_),
    .B1(_05718_),
    .X(_05726_));
 sky130_fd_sc_hd__o311a_1 _16366_ (.A1(net301),
    .A2(net300),
    .A3(_05699_),
    .B1(net386),
    .C1(_05717_),
    .X(_05727_));
 sky130_fd_sc_hd__o221ai_4 _16367_ (.A1(_05501_),
    .A2(_05523_),
    .B1(net275),
    .B2(_05699_),
    .C1(_05717_),
    .Y(_05728_));
 sky130_fd_sc_hd__o211ai_4 _16368_ (.A1(net398),
    .A2(net397),
    .B1(_05708_),
    .C1(_05710_),
    .Y(_05729_));
 sky130_fd_sc_hd__o221ai_4 _16369_ (.A1(_05465_),
    .A2(_05471_),
    .B1(net387),
    .B2(_05719_),
    .C1(_05728_),
    .Y(_05730_));
 sky130_fd_sc_hd__a21o_1 _16370_ (.A1(_05728_),
    .A2(_05729_),
    .B1(_05722_),
    .X(_05732_));
 sky130_fd_sc_hd__o211ai_2 _16371_ (.A1(net297),
    .A2(_05232_),
    .B1(_05730_),
    .C1(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__and3_2 _16372_ (.A(_05234_),
    .B(_05708_),
    .C(_05710_),
    .X(_05734_));
 sky130_fd_sc_hd__a31o_1 _16373_ (.A1(_05732_),
    .A2(net274),
    .A3(_05730_),
    .B1(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__nand3_1 _16374_ (.A(_05726_),
    .B(net403),
    .C(_05725_),
    .Y(_05736_));
 sky130_fd_sc_hd__a31o_1 _16375_ (.A1(_05732_),
    .A2(net274),
    .A3(_05730_),
    .B1(net403),
    .X(_05737_));
 sky130_fd_sc_hd__a311oi_4 _16376_ (.A1(_05732_),
    .A2(net274),
    .A3(_05730_),
    .B1(_05734_),
    .C1(net403),
    .Y(_05738_));
 sky130_fd_sc_hd__o221ai_4 _16377_ (.A1(_05196_),
    .A2(_05218_),
    .B1(net274),
    .B2(_05719_),
    .C1(_05733_),
    .Y(_05739_));
 sky130_fd_sc_hd__a31oi_2 _16378_ (.A1(_05726_),
    .A2(net403),
    .A3(_05725_),
    .B1(_05488_),
    .Y(_05740_));
 sky130_fd_sc_hd__a31o_2 _16379_ (.A1(_05726_),
    .A2(net403),
    .A3(_05725_),
    .B1(_05488_),
    .X(_05741_));
 sky130_fd_sc_hd__o2bb2ai_2 _16380_ (.A1_N(_05736_),
    .A2_N(_05739_),
    .B1(_03289_),
    .B2(_05476_),
    .Y(_05743_));
 sky130_fd_sc_hd__a31o_1 _16381_ (.A1(net403),
    .A2(_05725_),
    .A3(_05726_),
    .B1(_05489_),
    .X(_05744_));
 sky130_fd_sc_hd__o22a_1 _16382_ (.A1(_05481_),
    .A2(net269),
    .B1(_05738_),
    .B2(_05744_),
    .X(_05745_));
 sky130_fd_sc_hd__o211ai_1 _16383_ (.A1(_05738_),
    .A2(_05744_),
    .B1(_05485_),
    .C1(_05743_),
    .Y(_05746_));
 sky130_fd_sc_hd__o21ai_1 _16384_ (.A1(_05478_),
    .A2(_05479_),
    .B1(_05735_),
    .Y(_05747_));
 sky130_fd_sc_hd__a22oi_4 _16385_ (.A1(_05486_),
    .A2(_05735_),
    .B1(_05745_),
    .B2(_05743_),
    .Y(_05748_));
 sky130_fd_sc_hd__or4_4 _16386_ (.A(net36),
    .B(net37),
    .C(net38),
    .D(_03975_),
    .X(_05749_));
 sky130_fd_sc_hd__a21boi_4 _16387_ (.A1(_05749_),
    .A2(net409),
    .B1_N(net39),
    .Y(_05750_));
 sky130_fd_sc_hd__and3b_4 _16388_ (.A_N(net39),
    .B(_05749_),
    .C(net409),
    .X(_05751_));
 sky130_fd_sc_hd__or2_4 _16389_ (.A(net265),
    .B(net264),
    .X(_05752_));
 sky130_fd_sc_hd__nor2_8 _16390_ (.A(net265),
    .B(net264),
    .Y(_05754_));
 sky130_fd_sc_hd__o2bb2a_1 _16391_ (.A1_N(_05746_),
    .A2_N(_05747_),
    .B1(_05754_),
    .B2(_03289_),
    .X(_05755_));
 sky130_fd_sc_hd__a21oi_1 _16392_ (.A1(_05746_),
    .A2(_05747_),
    .B1(_03289_),
    .Y(_05756_));
 sky130_fd_sc_hd__a31oi_2 _16393_ (.A1(net1),
    .A2(_05748_),
    .A3(net241),
    .B1(_05755_),
    .Y(_05757_));
 sky130_fd_sc_hd__xnor2_1 _16394_ (.A(_05495_),
    .B(_05757_),
    .Y(net71));
 sky130_fd_sc_hd__nand3_1 _16395_ (.A(_05237_),
    .B(_05757_),
    .C(_05492_),
    .Y(_05758_));
 sky130_fd_sc_hd__or4_4 _16396_ (.A(net5),
    .B(net6),
    .C(net7),
    .D(_04150_),
    .X(_05759_));
 sky130_fd_sc_hd__and3b_4 _16397_ (.A_N(net8),
    .B(_05759_),
    .C(net410),
    .X(_05760_));
 sky130_fd_sc_hd__or3b_4 _16398_ (.A(_03399_),
    .B(net8),
    .C_N(_05759_),
    .X(_05761_));
 sky130_fd_sc_hd__a21boi_4 _16399_ (.A1(_05759_),
    .A2(net410),
    .B1_N(net8),
    .Y(_05762_));
 sky130_fd_sc_hd__a21bo_4 _16400_ (.A1(_05759_),
    .A2(net410),
    .B1_N(net8),
    .X(_05764_));
 sky130_fd_sc_hd__o311a_4 _16401_ (.A1(net6),
    .A2(net7),
    .A3(_05241_),
    .B1(net8),
    .C1(net410),
    .X(_05765_));
 sky130_fd_sc_hd__a21oi_4 _16402_ (.A1(_05759_),
    .A2(net410),
    .B1(net8),
    .Y(_05766_));
 sky130_fd_sc_hd__nor2_8 _16403_ (.A(_05760_),
    .B(_05762_),
    .Y(_05767_));
 sky130_fd_sc_hd__nor2_8 _16404_ (.A(_05765_),
    .B(_05766_),
    .Y(_05768_));
 sky130_fd_sc_hd__or3_1 _16405_ (.A(_03178_),
    .B(_05765_),
    .C(net289),
    .X(_05769_));
 sky130_fd_sc_hd__o221a_2 _16406_ (.A1(net408),
    .A2(_05152_),
    .B1(_05760_),
    .B2(net290),
    .C1(net33),
    .X(_05770_));
 sky130_fd_sc_hd__or4_1 _16407_ (.A(_03178_),
    .B(_05174_),
    .C(_05765_),
    .D(net289),
    .X(_05771_));
 sky130_fd_sc_hd__a22oi_2 _16408_ (.A1(net291),
    .A2(_05251_),
    .B1(_05515_),
    .B2(_05511_),
    .Y(_05772_));
 sky130_fd_sc_hd__o2bb2ai_1 _16409_ (.A1_N(_05511_),
    .A2_N(_05515_),
    .B1(_05252_),
    .B2(net267),
    .Y(_05773_));
 sky130_fd_sc_hd__a211o_1 _16410_ (.A1(net261),
    .A2(net33),
    .B1(_05500_),
    .C1(_05503_),
    .X(_05775_));
 sky130_fd_sc_hd__o31a_1 _16411_ (.A1(_05509_),
    .A2(_05765_),
    .A3(net289),
    .B1(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__o21ai_4 _16412_ (.A1(_05509_),
    .A2(net262),
    .B1(_05775_),
    .Y(_05777_));
 sky130_fd_sc_hd__nand2_2 _16413_ (.A(_05773_),
    .B(_05776_),
    .Y(_05778_));
 sky130_fd_sc_hd__o211ai_4 _16414_ (.A1(net267),
    .A2(_05252_),
    .B1(_05777_),
    .C1(_05517_),
    .Y(_05779_));
 sky130_fd_sc_hd__nand2_1 _16415_ (.A(_05778_),
    .B(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__nand3_1 _16416_ (.A(_05778_),
    .B(_05779_),
    .C(_05174_),
    .Y(_05781_));
 sky130_fd_sc_hd__o32a_2 _16417_ (.A1(_03178_),
    .A2(_05765_),
    .A3(net289),
    .B1(net408),
    .B2(_05152_),
    .X(_05782_));
 sky130_fd_sc_hd__a21oi_1 _16418_ (.A1(_05778_),
    .A2(_05779_),
    .B1(_05185_),
    .Y(_05783_));
 sky130_fd_sc_hd__a31o_2 _16419_ (.A1(_05778_),
    .A2(_05779_),
    .A3(_05174_),
    .B1(_05770_),
    .X(_05784_));
 sky130_fd_sc_hd__and3_1 _16420_ (.A(_05359_),
    .B(_05381_),
    .C(_05784_),
    .X(_05786_));
 sky130_fd_sc_hd__or4_2 _16421_ (.A(net402),
    .B(net400),
    .C(_05782_),
    .D(_05783_),
    .X(_05787_));
 sky130_fd_sc_hd__a311oi_4 _16422_ (.A1(_05778_),
    .A2(_05779_),
    .A3(_05174_),
    .B1(net293),
    .C1(_05770_),
    .Y(_05788_));
 sky130_fd_sc_hd__a311o_2 _16423_ (.A1(_05778_),
    .A2(_05779_),
    .A3(_05174_),
    .B1(net293),
    .C1(_05770_),
    .X(_05789_));
 sky130_fd_sc_hd__a22o_1 _16424_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_05780_),
    .B2(_05174_),
    .X(_05790_));
 sky130_fd_sc_hd__a21oi_2 _16425_ (.A1(_05771_),
    .A2(_05781_),
    .B1(net295),
    .Y(_05791_));
 sky130_fd_sc_hd__o21ai_4 _16426_ (.A1(_05242_),
    .A2(net317),
    .B1(_05784_),
    .Y(_05792_));
 sky130_fd_sc_hd__nand2_1 _16427_ (.A(_05789_),
    .B(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__a22oi_2 _16428_ (.A1(_05522_),
    .A2(_05529_),
    .B1(_05538_),
    .B2(_05528_),
    .Y(_05794_));
 sky130_fd_sc_hd__o22ai_2 _16429_ (.A1(_05521_),
    .A2(_05530_),
    .B1(_05527_),
    .B2(_05539_),
    .Y(_05795_));
 sky130_fd_sc_hd__o211ai_4 _16430_ (.A1(_05790_),
    .A2(_05782_),
    .B1(_05789_),
    .C1(_05795_),
    .Y(_05797_));
 sky130_fd_sc_hd__o221ai_4 _16431_ (.A1(net299),
    .A2(_05524_),
    .B1(_05788_),
    .B2(_05791_),
    .C1(_05541_),
    .Y(_05798_));
 sky130_fd_sc_hd__o211ai_2 _16432_ (.A1(net402),
    .A2(net400),
    .B1(_05797_),
    .C1(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__a211o_2 _16433_ (.A1(_05787_),
    .A2(_05799_),
    .B1(net384),
    .C1(net383),
    .X(_05800_));
 sky130_fd_sc_hd__a2bb2oi_2 _16434_ (.A1_N(net339),
    .A2_N(_04184_),
    .B1(_05787_),
    .B2(_05799_),
    .Y(_05801_));
 sky130_fd_sc_hd__a22o_1 _16435_ (.A1(_04173_),
    .A2(_04195_),
    .B1(_05787_),
    .B2(_05799_),
    .X(_05802_));
 sky130_fd_sc_hd__a311oi_4 _16436_ (.A1(net388),
    .A2(_05797_),
    .A3(_05798_),
    .B1(net298),
    .C1(_05786_),
    .Y(_05803_));
 sky130_fd_sc_hd__a311o_2 _16437_ (.A1(net388),
    .A2(_05797_),
    .A3(_05798_),
    .B1(net298),
    .C1(_05786_),
    .X(_05804_));
 sky130_fd_sc_hd__a31oi_2 _16438_ (.A1(_05297_),
    .A2(_05547_),
    .A3(_05553_),
    .B1(_05550_),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_2 _16439_ (.A1(_02137_),
    .A2(_05544_),
    .B1(_05559_),
    .Y(_05806_));
 sky130_fd_sc_hd__nand3_1 _16440_ (.A(_05802_),
    .B(_05804_),
    .C(_05806_),
    .Y(_05808_));
 sky130_fd_sc_hd__o21ai_1 _16441_ (.A1(_05801_),
    .A2(_05803_),
    .B1(_05805_),
    .Y(_05809_));
 sky130_fd_sc_hd__nand3_4 _16442_ (.A(_05809_),
    .B(net359),
    .C(_05808_),
    .Y(_05810_));
 sky130_fd_sc_hd__nand2_2 _16443_ (.A(_05800_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__a2bb2oi_2 _16444_ (.A1_N(_02049_),
    .A2_N(net342),
    .B1(_05800_),
    .B2(_05810_),
    .Y(_05812_));
 sky130_fd_sc_hd__a22o_2 _16445_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_05800_),
    .B2(_05810_),
    .X(_05813_));
 sky130_fd_sc_hd__and3_1 _16446_ (.A(_05810_),
    .B(_02137_),
    .C(_05800_),
    .X(_05814_));
 sky130_fd_sc_hd__nand3_2 _16447_ (.A(_05810_),
    .B(_02137_),
    .C(_05800_),
    .Y(_05815_));
 sky130_fd_sc_hd__o2111a_2 _16448_ (.A1(_02729_),
    .A2(_02510_),
    .B1(_02696_),
    .C1(_04855_),
    .D1(_04877_),
    .X(_05816_));
 sky130_fd_sc_hd__o2111ai_1 _16449_ (.A1(_02729_),
    .A2(_02510_),
    .B1(_02696_),
    .C1(_04855_),
    .D1(_04877_),
    .Y(_05817_));
 sky130_fd_sc_hd__nor3_1 _16450_ (.A(_05817_),
    .B(_05314_),
    .C(_05312_),
    .Y(_05819_));
 sky130_fd_sc_hd__nand4_4 _16451_ (.A(_05313_),
    .B(_05315_),
    .C(_05816_),
    .D(_02707_),
    .Y(_05820_));
 sky130_fd_sc_hd__nand4_2 _16452_ (.A(_05816_),
    .B(_05569_),
    .C(_05315_),
    .D(_05313_),
    .Y(_05821_));
 sky130_fd_sc_hd__nor2_1 _16453_ (.A(_05570_),
    .B(_05820_),
    .Y(_05822_));
 sky130_fd_sc_hd__nand4_2 _16454_ (.A(_05566_),
    .B(_05819_),
    .C(_05569_),
    .D(_02707_),
    .Y(_05823_));
 sky130_fd_sc_hd__a41oi_4 _16455_ (.A1(_05816_),
    .A2(_05569_),
    .A3(_05315_),
    .A4(_05313_),
    .B1(_05565_),
    .Y(_05824_));
 sky130_fd_sc_hd__o211a_1 _16456_ (.A1(_05572_),
    .A2(_05568_),
    .B1(_05566_),
    .C1(_05821_),
    .X(_05825_));
 sky130_fd_sc_hd__o211ai_4 _16457_ (.A1(_05568_),
    .A2(_05572_),
    .B1(_05821_),
    .C1(_05566_),
    .Y(_05826_));
 sky130_fd_sc_hd__a2bb2oi_4 _16458_ (.A1_N(_05570_),
    .A2_N(_05820_),
    .B1(_05576_),
    .B2(_05824_),
    .Y(_05827_));
 sky130_fd_sc_hd__o21a_1 _16459_ (.A1(_05570_),
    .A2(_05820_),
    .B1(_05815_),
    .X(_05828_));
 sky130_fd_sc_hd__o21ai_1 _16460_ (.A1(_05570_),
    .A2(_05820_),
    .B1(_05815_),
    .Y(_05830_));
 sky130_fd_sc_hd__a41oi_2 _16461_ (.A1(_02060_),
    .A2(_02082_),
    .A3(_05800_),
    .A4(_05810_),
    .B1(_05812_),
    .Y(_05831_));
 sky130_fd_sc_hd__nor3_1 _16462_ (.A(_05812_),
    .B(_05830_),
    .C(_05825_),
    .Y(_05832_));
 sky130_fd_sc_hd__nand4_4 _16463_ (.A(_05813_),
    .B(_05815_),
    .C(_05823_),
    .D(_05826_),
    .Y(_05833_));
 sky130_fd_sc_hd__o22ai_4 _16464_ (.A1(_05812_),
    .A2(_05814_),
    .B1(_05822_),
    .B2(_05825_),
    .Y(_05834_));
 sky130_fd_sc_hd__o22ai_2 _16465_ (.A1(net379),
    .A2(net378),
    .B1(_05827_),
    .B2(_05831_),
    .Y(_05835_));
 sky130_fd_sc_hd__nand3_2 _16466_ (.A(_05834_),
    .B(net357),
    .C(_05833_),
    .Y(_05836_));
 sky130_fd_sc_hd__and3_4 _16467_ (.A(_06804_),
    .B(_06826_),
    .C(_05811_),
    .X(_05837_));
 sky130_fd_sc_hd__a211o_2 _16468_ (.A1(_05800_),
    .A2(_05810_),
    .B1(net379),
    .C1(net378),
    .X(_05838_));
 sky130_fd_sc_hd__a31oi_4 _16469_ (.A1(_05834_),
    .A2(net357),
    .A3(_05833_),
    .B1(_05837_),
    .Y(_05839_));
 sky130_fd_sc_hd__a21oi_2 _16470_ (.A1(_05836_),
    .A2(_05838_),
    .B1(net356),
    .Y(_05841_));
 sky130_fd_sc_hd__or3_2 _16471_ (.A(net372),
    .B(net371),
    .C(_05839_),
    .X(_05842_));
 sky130_fd_sc_hd__o22ai_4 _16472_ (.A1(_00218_),
    .A2(_00229_),
    .B1(_05832_),
    .B2(_05835_),
    .Y(_05843_));
 sky130_fd_sc_hd__a311oi_4 _16473_ (.A1(_05834_),
    .A2(net357),
    .A3(_05833_),
    .B1(_05837_),
    .C1(net319),
    .Y(_05844_));
 sky130_fd_sc_hd__a31o_1 _16474_ (.A1(_06804_),
    .A2(_06826_),
    .A3(_05811_),
    .B1(_05843_),
    .X(_05845_));
 sky130_fd_sc_hd__a21oi_4 _16475_ (.A1(_05836_),
    .A2(_05838_),
    .B1(net320),
    .Y(_05846_));
 sky130_fd_sc_hd__a21o_1 _16476_ (.A1(_05836_),
    .A2(_05838_),
    .B1(net320),
    .X(_05847_));
 sky130_fd_sc_hd__a31o_2 _16477_ (.A1(_05330_),
    .A2(_05583_),
    .A3(_05586_),
    .B1(_05587_),
    .X(_05848_));
 sky130_fd_sc_hd__a31oi_4 _16478_ (.A1(_05330_),
    .A2(_05583_),
    .A3(_05586_),
    .B1(_05587_),
    .Y(_05849_));
 sky130_fd_sc_hd__o21ai_4 _16479_ (.A1(_05844_),
    .A2(_05846_),
    .B1(_05849_),
    .Y(_05850_));
 sky130_fd_sc_hd__o211ai_4 _16480_ (.A1(_05837_),
    .A2(_05843_),
    .B1(_05848_),
    .C1(_05847_),
    .Y(_05852_));
 sky130_fd_sc_hd__nand3_4 _16481_ (.A(_05850_),
    .B(_05852_),
    .C(net356),
    .Y(_05853_));
 sky130_fd_sc_hd__a31oi_4 _16482_ (.A1(_05850_),
    .A2(_05852_),
    .A3(net356),
    .B1(_05841_),
    .Y(_05854_));
 sky130_fd_sc_hd__inv_2 _16483_ (.A(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__o221a_1 _16484_ (.A1(_05349_),
    .A2(_05350_),
    .B1(net331),
    .B2(_05598_),
    .C1(_05346_),
    .X(_05856_));
 sky130_fd_sc_hd__o31a_1 _16485_ (.A1(_11210_),
    .A2(_11232_),
    .A3(_05597_),
    .B1(_05606_),
    .X(_05857_));
 sky130_fd_sc_hd__o21ai_1 _16486_ (.A1(_05607_),
    .A2(_05603_),
    .B1(_05601_),
    .Y(_05858_));
 sky130_fd_sc_hd__o2bb2ai_2 _16487_ (.A1_N(_05601_),
    .A2_N(_05607_),
    .B1(_05602_),
    .B2(_05593_),
    .Y(_05859_));
 sky130_fd_sc_hd__a31oi_1 _16488_ (.A1(_05850_),
    .A2(_05852_),
    .A3(net356),
    .B1(net325),
    .Y(_05860_));
 sky130_fd_sc_hd__a311oi_4 _16489_ (.A1(_05850_),
    .A2(_05852_),
    .A3(net356),
    .B1(net325),
    .C1(_05841_),
    .Y(_05861_));
 sky130_fd_sc_hd__o221ai_4 _16490_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_05839_),
    .B2(net356),
    .C1(_05853_),
    .Y(_05863_));
 sky130_fd_sc_hd__a2bb2oi_4 _16491_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_05842_),
    .B2(_05853_),
    .Y(_05864_));
 sky130_fd_sc_hd__a2bb2o_1 _16492_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_05842_),
    .B2(_05853_),
    .X(_05865_));
 sky130_fd_sc_hd__o211ai_1 _16493_ (.A1(_05603_),
    .A2(_05856_),
    .B1(_05863_),
    .C1(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__o22ai_1 _16494_ (.A1(_05599_),
    .A2(_05857_),
    .B1(_05861_),
    .B2(_05864_),
    .Y(_05867_));
 sky130_fd_sc_hd__o21ai_1 _16495_ (.A1(_12888_),
    .A2(_05854_),
    .B1(_05858_),
    .Y(_05868_));
 sky130_fd_sc_hd__o22ai_2 _16496_ (.A1(_05603_),
    .A2(_05856_),
    .B1(_05861_),
    .B2(_05864_),
    .Y(_05869_));
 sky130_fd_sc_hd__nand3_1 _16497_ (.A(_05866_),
    .B(_05867_),
    .C(_08721_),
    .Y(_05870_));
 sky130_fd_sc_hd__or3_1 _16498_ (.A(net353),
    .B(net352),
    .C(_05854_),
    .X(_05871_));
 sky130_fd_sc_hd__o221ai_4 _16499_ (.A1(net353),
    .A2(net352),
    .B1(_05861_),
    .B2(_05868_),
    .C1(_05869_),
    .Y(_05872_));
 sky130_fd_sc_hd__o21ai_2 _16500_ (.A1(_08721_),
    .A2(_05854_),
    .B1(_05872_),
    .Y(_05874_));
 sky130_fd_sc_hd__o211ai_4 _16501_ (.A1(_08721_),
    .A2(_05854_),
    .B1(net331),
    .C1(_05872_),
    .Y(_05875_));
 sky130_fd_sc_hd__a2bb2oi_1 _16502_ (.A1_N(_11210_),
    .A2_N(_11232_),
    .B1(_05871_),
    .B2(_05872_),
    .Y(_05876_));
 sky130_fd_sc_hd__o211ai_4 _16503_ (.A1(_05855_),
    .A2(_08721_),
    .B1(net330),
    .C1(_05870_),
    .Y(_05877_));
 sky130_fd_sc_hd__o221a_1 _16504_ (.A1(_08907_),
    .A2(_05362_),
    .B1(_10015_),
    .B2(_05616_),
    .C1(_05623_),
    .X(_05878_));
 sky130_fd_sc_hd__a21oi_2 _16505_ (.A1(_05619_),
    .A2(_05625_),
    .B1(_05620_),
    .Y(_05879_));
 sky130_fd_sc_hd__o21ai_1 _16506_ (.A1(_05618_),
    .A2(_05624_),
    .B1(_05621_),
    .Y(_05880_));
 sky130_fd_sc_hd__o2bb2ai_4 _16507_ (.A1_N(_05875_),
    .A2_N(_05877_),
    .B1(_05878_),
    .B2(_05620_),
    .Y(_05881_));
 sky130_fd_sc_hd__nand3_4 _16508_ (.A(_05875_),
    .B(_05877_),
    .C(_05879_),
    .Y(_05882_));
 sky130_fd_sc_hd__nand3_2 _16509_ (.A(_05881_),
    .B(_05882_),
    .C(net337),
    .Y(_05883_));
 sky130_fd_sc_hd__and3_2 _16510_ (.A(_05874_),
    .B(_09818_),
    .C(_09796_),
    .X(_05885_));
 sky130_fd_sc_hd__a211o_1 _16511_ (.A1(_05871_),
    .A2(_05872_),
    .B1(net350),
    .C1(net349),
    .X(_05886_));
 sky130_fd_sc_hd__a31oi_4 _16512_ (.A1(_05881_),
    .A2(_05882_),
    .A3(net337),
    .B1(_05885_),
    .Y(_05887_));
 sky130_fd_sc_hd__a22oi_4 _16513_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_05883_),
    .B2(_05886_),
    .Y(_05888_));
 sky130_fd_sc_hd__a22o_1 _16514_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_05883_),
    .B2(_05886_),
    .X(_05889_));
 sky130_fd_sc_hd__a21oi_4 _16515_ (.A1(_05638_),
    .A2(_05640_),
    .B1(_05641_),
    .Y(_05890_));
 sky130_fd_sc_hd__a32o_2 _16516_ (.A1(_08918_),
    .A2(_05617_),
    .A3(_05630_),
    .B1(_05638_),
    .B2(_05640_),
    .X(_05891_));
 sky130_fd_sc_hd__a311oi_4 _16517_ (.A1(_05881_),
    .A2(_05882_),
    .A3(net337),
    .B1(net348),
    .C1(_05885_),
    .Y(_05892_));
 sky130_fd_sc_hd__a311o_2 _16518_ (.A1(_05881_),
    .A2(_05882_),
    .A3(net337),
    .B1(net348),
    .C1(_05885_),
    .X(_05893_));
 sky130_fd_sc_hd__nand3_2 _16519_ (.A(_05889_),
    .B(_05891_),
    .C(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__o21ai_2 _16520_ (.A1(_05888_),
    .A2(_05892_),
    .B1(_05890_),
    .Y(_05896_));
 sky130_fd_sc_hd__o211ai_4 _16521_ (.A1(net347),
    .A2(net346),
    .B1(_05894_),
    .C1(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__a21oi_1 _16522_ (.A1(_05883_),
    .A2(_05886_),
    .B1(net334),
    .Y(_05898_));
 sky130_fd_sc_hd__or3_2 _16523_ (.A(net347),
    .B(net346),
    .C(_05887_),
    .X(_05899_));
 sky130_fd_sc_hd__a31oi_4 _16524_ (.A1(_05896_),
    .A2(net334),
    .A3(_05894_),
    .B1(_05898_),
    .Y(_05900_));
 sky130_fd_sc_hd__o221ai_4 _16525_ (.A1(_05238_),
    .A2(_05396_),
    .B1(_05647_),
    .B2(_07888_),
    .C1(_05399_),
    .Y(_05901_));
 sky130_fd_sc_hd__a31o_1 _16526_ (.A1(_05397_),
    .A2(_05650_),
    .A3(_05653_),
    .B1(_05655_),
    .X(_05902_));
 sky130_fd_sc_hd__o211ai_4 _16527_ (.A1(_07888_),
    .A2(_05647_),
    .B1(_08907_),
    .C1(_05657_),
    .Y(_05903_));
 sky130_fd_sc_hd__o211ai_4 _16528_ (.A1(_08819_),
    .A2(net367),
    .B1(_05653_),
    .C1(_05901_),
    .Y(_05904_));
 sky130_fd_sc_hd__and4_2 _16529_ (.A(_05904_),
    .B(net313),
    .C(_05903_),
    .D(_05900_),
    .X(_05905_));
 sky130_fd_sc_hd__nand4_1 _16530_ (.A(_05904_),
    .B(_05900_),
    .C(net313),
    .D(_05903_),
    .Y(_05907_));
 sky130_fd_sc_hd__a31oi_4 _16531_ (.A1(_05904_),
    .A2(net313),
    .A3(_05903_),
    .B1(_05900_),
    .Y(_05908_));
 sky130_fd_sc_hd__a31o_1 _16532_ (.A1(_05904_),
    .A2(net313),
    .A3(_05903_),
    .B1(_05900_),
    .X(_05909_));
 sky130_fd_sc_hd__o211ai_2 _16533_ (.A1(net334),
    .A2(_05887_),
    .B1(_08907_),
    .C1(_05897_),
    .Y(_05910_));
 sky130_fd_sc_hd__a22oi_4 _16534_ (.A1(_08830_),
    .A2(_08852_),
    .B1(_05897_),
    .B2(_05899_),
    .Y(_05911_));
 sky130_fd_sc_hd__o22a_2 _16535_ (.A1(_14458_),
    .A2(_00000_),
    .B1(_05905_),
    .B2(_05908_),
    .X(_05912_));
 sky130_fd_sc_hd__a211o_2 _16536_ (.A1(_05907_),
    .A2(_05909_),
    .B1(net324),
    .C1(net322),
    .X(_05913_));
 sky130_fd_sc_hd__o221a_1 _16537_ (.A1(_05418_),
    .A2(_05415_),
    .B1(_07033_),
    .B2(_05662_),
    .C1(_05413_),
    .X(_05914_));
 sky130_fd_sc_hd__o21ai_2 _16538_ (.A1(_07033_),
    .A2(_05662_),
    .B1(_05496_),
    .Y(_05915_));
 sky130_fd_sc_hd__o32a_1 _16539_ (.A1(_06945_),
    .A2(net377),
    .A3(_05663_),
    .B1(_05668_),
    .B2(_05497_),
    .X(_05916_));
 sky130_fd_sc_hd__nor3_4 _16540_ (.A(_05908_),
    .B(_07899_),
    .C(_05905_),
    .Y(_05918_));
 sky130_fd_sc_hd__nand3_2 _16541_ (.A(_05909_),
    .B(_07888_),
    .C(_05907_),
    .Y(_05919_));
 sky130_fd_sc_hd__o22a_2 _16542_ (.A1(net389),
    .A2(net370),
    .B1(_05905_),
    .B2(_05908_),
    .X(_05920_));
 sky130_fd_sc_hd__o22ai_4 _16543_ (.A1(net389),
    .A2(net370),
    .B1(_05905_),
    .B2(_05908_),
    .Y(_05921_));
 sky130_fd_sc_hd__o211ai_4 _16544_ (.A1(_07044_),
    .A2(_05663_),
    .B1(_05915_),
    .C1(_05919_),
    .Y(_05922_));
 sky130_fd_sc_hd__o2111ai_4 _16545_ (.A1(_07044_),
    .A2(_05663_),
    .B1(_05915_),
    .C1(_05919_),
    .D1(_05921_),
    .Y(_05923_));
 sky130_fd_sc_hd__o22ai_4 _16546_ (.A1(_05667_),
    .A2(_05914_),
    .B1(_05918_),
    .B2(_05920_),
    .Y(_05924_));
 sky130_fd_sc_hd__o211ai_4 _16547_ (.A1(_05920_),
    .A2(_05922_),
    .B1(net310),
    .C1(_05924_),
    .Y(_05925_));
 sky130_fd_sc_hd__a31oi_4 _16548_ (.A1(_05924_),
    .A2(net310),
    .A3(_05923_),
    .B1(_05912_),
    .Y(_05926_));
 sky130_fd_sc_hd__and3_2 _16549_ (.A(_01973_),
    .B(_05913_),
    .C(_05925_),
    .X(_05927_));
 sky130_fd_sc_hd__a21oi_2 _16550_ (.A1(_05686_),
    .A2(_05689_),
    .B1(_05683_),
    .Y(_05929_));
 sky130_fd_sc_hd__a311oi_4 _16551_ (.A1(_05924_),
    .A2(net310),
    .A3(_05923_),
    .B1(_05912_),
    .C1(_07044_),
    .Y(_05930_));
 sky130_fd_sc_hd__a311o_1 _16552_ (.A1(_05924_),
    .A2(net310),
    .A3(_05923_),
    .B1(_05912_),
    .C1(_07044_),
    .X(_05931_));
 sky130_fd_sc_hd__a2bb2oi_4 _16553_ (.A1_N(_06945_),
    .A2_N(net377),
    .B1(_05913_),
    .B2(_05925_),
    .Y(_05932_));
 sky130_fd_sc_hd__a22o_1 _16554_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_05913_),
    .B2(_05925_),
    .X(_05933_));
 sky130_fd_sc_hd__o2bb2ai_1 _16555_ (.A1_N(_05684_),
    .A2_N(_05693_),
    .B1(_05926_),
    .B2(_07033_),
    .Y(_05934_));
 sky130_fd_sc_hd__nand3b_2 _16556_ (.A_N(_05929_),
    .B(_05931_),
    .C(_05933_),
    .Y(_05935_));
 sky130_fd_sc_hd__o21ai_4 _16557_ (.A1(_05930_),
    .A2(_05932_),
    .B1(_05929_),
    .Y(_05936_));
 sky130_fd_sc_hd__a21oi_4 _16558_ (.A1(_05935_),
    .A2(_05936_),
    .B1(_01973_),
    .Y(_05937_));
 sky130_fd_sc_hd__or3_2 _16559_ (.A(net305),
    .B(net303),
    .C(_05926_),
    .X(_05938_));
 sky130_fd_sc_hd__o221ai_4 _16560_ (.A1(net305),
    .A2(net303),
    .B1(_05930_),
    .B2(_05934_),
    .C1(_05936_),
    .Y(_05940_));
 sky130_fd_sc_hd__a21oi_2 _16561_ (.A1(_05938_),
    .A2(_05940_),
    .B1(net275),
    .Y(_05941_));
 sky130_fd_sc_hd__o21ai_2 _16562_ (.A1(_05703_),
    .A2(_05713_),
    .B1(_05712_),
    .Y(_05942_));
 sky130_fd_sc_hd__a22oi_2 _16563_ (.A1(_05682_),
    .A2(_05711_),
    .B1(_05702_),
    .B2(_05714_),
    .Y(_05943_));
 sky130_fd_sc_hd__a2bb2oi_4 _16564_ (.A1_N(_06245_),
    .A2_N(_06267_),
    .B1(_05938_),
    .B2(_05940_),
    .Y(_05944_));
 sky130_fd_sc_hd__a31oi_1 _16565_ (.A1(_05935_),
    .A2(_05936_),
    .A3(_01962_),
    .B1(_06343_),
    .Y(_05945_));
 sky130_fd_sc_hd__o221a_2 _16566_ (.A1(_06289_),
    .A2(net391),
    .B1(_01962_),
    .B2(_05926_),
    .C1(_05940_),
    .X(_05946_));
 sky130_fd_sc_hd__o221ai_4 _16567_ (.A1(_06289_),
    .A2(net391),
    .B1(_01962_),
    .B2(_05926_),
    .C1(_05940_),
    .Y(_05947_));
 sky130_fd_sc_hd__nand2_1 _16568_ (.A(_05943_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__a211oi_1 _16569_ (.A1(_05945_),
    .A2(_05938_),
    .B1(_05942_),
    .C1(_05944_),
    .Y(_05949_));
 sky130_fd_sc_hd__o21a_1 _16570_ (.A1(_05944_),
    .A2(_05946_),
    .B1(_05942_),
    .X(_05951_));
 sky130_fd_sc_hd__o21ai_1 _16571_ (.A1(_05944_),
    .A2(_05946_),
    .B1(_05942_),
    .Y(_05952_));
 sky130_fd_sc_hd__o211a_1 _16572_ (.A1(_05944_),
    .A2(_05948_),
    .B1(net275),
    .C1(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__o211ai_2 _16573_ (.A1(_05944_),
    .A2(_05948_),
    .B1(net275),
    .C1(_05952_),
    .Y(_05954_));
 sky130_fd_sc_hd__o22ai_1 _16574_ (.A1(net301),
    .A2(net300),
    .B1(_05949_),
    .B2(_05951_),
    .Y(_05955_));
 sky130_fd_sc_hd__o21ai_1 _16575_ (.A1(_05927_),
    .A2(_05937_),
    .B1(_04040_),
    .Y(_05956_));
 sky130_fd_sc_hd__o31ai_4 _16576_ (.A1(net275),
    .A2(_05927_),
    .A3(_05937_),
    .B1(_05954_),
    .Y(_05957_));
 sky130_fd_sc_hd__o21ai_4 _16577_ (.A1(_05465_),
    .A2(_05471_),
    .B1(_05728_),
    .Y(_05958_));
 sky130_fd_sc_hd__o32ai_1 _16578_ (.A1(_05501_),
    .A2(_05523_),
    .A3(_05719_),
    .B1(_05721_),
    .B2(_05727_),
    .Y(_05959_));
 sky130_fd_sc_hd__o211ai_4 _16579_ (.A1(_05719_),
    .A2(net387),
    .B1(_05851_),
    .C1(_05958_),
    .Y(_05960_));
 sky130_fd_sc_hd__inv_2 _16580_ (.A(_05960_),
    .Y(_05962_));
 sky130_fd_sc_hd__a22oi_4 _16581_ (.A1(_05774_),
    .A2(_05796_),
    .B1(_05958_),
    .B2(_05729_),
    .Y(_05963_));
 sky130_fd_sc_hd__o2bb2ai_4 _16582_ (.A1_N(_05729_),
    .A2_N(_05958_),
    .B1(_05763_),
    .B2(_05785_),
    .Y(_05964_));
 sky130_fd_sc_hd__o2111a_1 _16583_ (.A1(_05941_),
    .A2(_05953_),
    .B1(net274),
    .C1(_05960_),
    .D1(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__o2111ai_4 _16584_ (.A1(_05941_),
    .A2(_05953_),
    .B1(net274),
    .C1(_05960_),
    .D1(_05964_),
    .Y(_05966_));
 sky130_fd_sc_hd__a31oi_1 _16585_ (.A1(_05964_),
    .A2(net274),
    .A3(_05960_),
    .B1(_05957_),
    .Y(_05967_));
 sky130_fd_sc_hd__a31o_2 _16586_ (.A1(_05964_),
    .A2(net274),
    .A3(_05960_),
    .B1(_05957_),
    .X(_05968_));
 sky130_fd_sc_hd__nor2_2 _16587_ (.A(_05965_),
    .B(_05967_),
    .Y(_05969_));
 sky130_fd_sc_hd__o2bb2ai_2 _16588_ (.A1_N(_05489_),
    .A2_N(_05736_),
    .B1(_05734_),
    .B2(_05737_),
    .Y(_05970_));
 sky130_fd_sc_hd__o22ai_4 _16589_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_05738_),
    .B2(_05740_),
    .Y(_05971_));
 sky130_fd_sc_hd__o211ai_4 _16590_ (.A1(net398),
    .A2(net397),
    .B1(_05739_),
    .C1(_05741_),
    .Y(_05973_));
 sky130_fd_sc_hd__o2111a_1 _16591_ (.A1(_05481_),
    .A2(net269),
    .B1(_05969_),
    .C1(_05971_),
    .D1(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__o2111ai_4 _16592_ (.A1(_05481_),
    .A2(net269),
    .B1(_05969_),
    .C1(_05971_),
    .D1(_05973_),
    .Y(_05975_));
 sky130_fd_sc_hd__a31oi_2 _16593_ (.A1(_05971_),
    .A2(_05973_),
    .A3(_05485_),
    .B1(_05969_),
    .Y(_05976_));
 sky130_fd_sc_hd__a31o_1 _16594_ (.A1(_05971_),
    .A2(_05973_),
    .A3(_05485_),
    .B1(_05969_),
    .X(_05977_));
 sky130_fd_sc_hd__o2111ai_4 _16595_ (.A1(_03399_),
    .A2(_05491_),
    .B1(_05534_),
    .C1(_05966_),
    .D1(_05968_),
    .Y(_05978_));
 sky130_fd_sc_hd__nor2_1 _16596_ (.A(_05974_),
    .B(_05976_),
    .Y(_05979_));
 sky130_fd_sc_hd__nand3_1 _16597_ (.A(_05977_),
    .B(net403),
    .C(_05975_),
    .Y(_05980_));
 sky130_fd_sc_hd__a21oi_2 _16598_ (.A1(_05975_),
    .A2(_05977_),
    .B1(net403),
    .Y(_05981_));
 sky130_fd_sc_hd__o21ai_2 _16599_ (.A1(_05974_),
    .A2(_05976_),
    .B1(_05250_),
    .Y(_05982_));
 sky130_fd_sc_hd__a21bo_1 _16600_ (.A1(_05980_),
    .A2(_05982_),
    .B1_N(_05756_),
    .X(_05984_));
 sky130_fd_sc_hd__a31oi_2 _16601_ (.A1(_05977_),
    .A2(net403),
    .A3(_05975_),
    .B1(_05756_),
    .Y(_05985_));
 sky130_fd_sc_hd__o21ai_4 _16602_ (.A1(_03289_),
    .A2(_05748_),
    .B1(_05980_),
    .Y(_05986_));
 sky130_fd_sc_hd__o211ai_4 _16603_ (.A1(_05981_),
    .A2(_05986_),
    .B1(net241),
    .C1(_05984_),
    .Y(_05987_));
 sky130_fd_sc_hd__o21ai_2 _16604_ (.A1(net241),
    .A2(_05979_),
    .B1(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__or4_4 _16605_ (.A(net37),
    .B(net38),
    .C(net39),
    .D(_05227_),
    .X(_05989_));
 sky130_fd_sc_hd__and3b_4 _16606_ (.A_N(net40),
    .B(_05989_),
    .C(net409),
    .X(_05990_));
 sky130_fd_sc_hd__nand3b_4 _16607_ (.A_N(net40),
    .B(_05989_),
    .C(net409),
    .Y(_05991_));
 sky130_fd_sc_hd__a21boi_4 _16608_ (.A1(_05989_),
    .A2(net409),
    .B1_N(net40),
    .Y(_05992_));
 sky130_fd_sc_hd__a21bo_4 _16609_ (.A1(_05989_),
    .A2(net409),
    .B1_N(net40),
    .X(_05993_));
 sky130_fd_sc_hd__nor2_8 _16610_ (.A(_05990_),
    .B(_05992_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand2_8 _16611_ (.A(_05991_),
    .B(_05993_),
    .Y(_05996_));
 sky130_fd_sc_hd__o221a_1 _16612_ (.A1(net241),
    .A2(_05979_),
    .B1(_05995_),
    .B2(_03289_),
    .C1(_05987_),
    .X(_05997_));
 sky130_fd_sc_hd__o311a_1 _16613_ (.A1(net266),
    .A2(_05751_),
    .A3(_05979_),
    .B1(net1),
    .C1(_05987_),
    .X(_05998_));
 sky130_fd_sc_hd__o211ai_1 _16614_ (.A1(net241),
    .A2(_05979_),
    .B1(net1),
    .C1(_05987_),
    .Y(_05999_));
 sky130_fd_sc_hd__a31o_1 _16615_ (.A1(net1),
    .A2(_05988_),
    .A3(_05996_),
    .B1(_05997_),
    .X(_06000_));
 sky130_fd_sc_hd__and3_1 _16616_ (.A(_05119_),
    .B(_05758_),
    .C(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__a21oi_1 _16617_ (.A1(_05119_),
    .A2(_05758_),
    .B1(_06000_),
    .Y(_06002_));
 sky130_fd_sc_hd__nor2_1 _16618_ (.A(_06001_),
    .B(_06002_),
    .Y(net72));
 sky130_fd_sc_hd__or2_1 _16619_ (.A(_05758_),
    .B(_06000_),
    .X(_06003_));
 sky130_fd_sc_hd__o211a_1 _16620_ (.A1(_05496_),
    .A2(_05667_),
    .B1(_05669_),
    .C1(_05921_),
    .X(_06005_));
 sky130_fd_sc_hd__nand2_1 _16621_ (.A(_05921_),
    .B(_05922_),
    .Y(_06006_));
 sky130_fd_sc_hd__a21oi_1 _16622_ (.A1(_05916_),
    .A2(_05919_),
    .B1(_05920_),
    .Y(_06007_));
 sky130_fd_sc_hd__or4_4 _16623_ (.A(net6),
    .B(net7),
    .C(net8),
    .D(_05241_),
    .X(_06008_));
 sky130_fd_sc_hd__and3b_4 _16624_ (.A_N(net9),
    .B(_06008_),
    .C(net410),
    .X(_06009_));
 sky130_fd_sc_hd__a21boi_4 _16625_ (.A1(_06008_),
    .A2(net410),
    .B1_N(net9),
    .Y(_06010_));
 sky130_fd_sc_hd__a21oi_4 _16626_ (.A1(_06008_),
    .A2(net410),
    .B1(net9),
    .Y(_06011_));
 sky130_fd_sc_hd__o311a_4 _16627_ (.A1(net7),
    .A2(net8),
    .A3(_05498_),
    .B1(net9),
    .C1(net410),
    .X(_06012_));
 sky130_fd_sc_hd__nor2_4 _16628_ (.A(_06009_),
    .B(net287),
    .Y(_06013_));
 sky130_fd_sc_hd__nor2_8 _16629_ (.A(net285),
    .B(_06012_),
    .Y(_06014_));
 sky130_fd_sc_hd__o21a_1 _16630_ (.A1(_06009_),
    .A2(_06010_),
    .B1(net33),
    .X(_06016_));
 sky130_fd_sc_hd__or3_4 _16631_ (.A(_03178_),
    .B(net286),
    .C(_06012_),
    .X(_06017_));
 sky130_fd_sc_hd__or4_2 _16632_ (.A(_03178_),
    .B(_05174_),
    .C(net286),
    .D(_06012_),
    .X(_06018_));
 sky130_fd_sc_hd__nor4_2 _16633_ (.A(_04327_),
    .B(_05257_),
    .C(_05514_),
    .D(_05777_),
    .Y(_06019_));
 sky130_fd_sc_hd__nand2_1 _16634_ (.A(_06019_),
    .B(_04404_),
    .Y(_06020_));
 sky130_fd_sc_hd__a31o_1 _16635_ (.A1(net33),
    .A2(net291),
    .A3(net261),
    .B1(_06019_),
    .X(_06021_));
 sky130_fd_sc_hd__a21oi_1 _16636_ (.A1(_05773_),
    .A2(_05776_),
    .B1(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__o21bai_4 _16637_ (.A1(_05777_),
    .A2(_05772_),
    .B1_N(_06021_),
    .Y(_06023_));
 sky130_fd_sc_hd__and3_2 _16638_ (.A(net261),
    .B(net253),
    .C(net33),
    .X(_06024_));
 sky130_fd_sc_hd__or4_2 _16639_ (.A(net286),
    .B(_03178_),
    .C(net262),
    .D(_06012_),
    .X(_06025_));
 sky130_fd_sc_hd__o32a_2 _16640_ (.A1(_03178_),
    .A2(net286),
    .A3(_06012_),
    .B1(_05765_),
    .B2(net289),
    .X(_06027_));
 sky130_fd_sc_hd__o2bb2ai_2 _16641_ (.A1_N(_06020_),
    .A2_N(_06023_),
    .B1(_06024_),
    .B2(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__a211oi_4 _16642_ (.A1(_06019_),
    .A2(_04404_),
    .B1(_06027_),
    .C1(_06024_),
    .Y(_06029_));
 sky130_fd_sc_hd__inv_2 _16643_ (.A(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__nand2_4 _16644_ (.A(_06023_),
    .B(_06029_),
    .Y(_06031_));
 sky130_fd_sc_hd__a21oi_1 _16645_ (.A1(_06023_),
    .A2(_06029_),
    .B1(_05185_),
    .Y(_06032_));
 sky130_fd_sc_hd__nand3_2 _16646_ (.A(_06028_),
    .B(_06031_),
    .C(_05174_),
    .Y(_06033_));
 sky130_fd_sc_hd__a21oi_2 _16647_ (.A1(_06028_),
    .A2(_06031_),
    .B1(_05185_),
    .Y(_06034_));
 sky130_fd_sc_hd__o31a_1 _16648_ (.A1(_03178_),
    .A2(_05174_),
    .A3(net254),
    .B1(_06033_),
    .X(_06035_));
 sky130_fd_sc_hd__o2bb2ai_2 _16649_ (.A1_N(_06032_),
    .A2_N(_06028_),
    .B1(_06017_),
    .B2(_05174_),
    .Y(_06036_));
 sky130_fd_sc_hd__and3_1 _16650_ (.A(_05359_),
    .B(_05381_),
    .C(_06036_),
    .X(_06038_));
 sky130_fd_sc_hd__a211o_2 _16651_ (.A1(_05185_),
    .A2(_06017_),
    .B1(net388),
    .C1(_06034_),
    .X(_06039_));
 sky130_fd_sc_hd__nand3_4 _16652_ (.A(_06033_),
    .B(net267),
    .C(_06018_),
    .Y(_06040_));
 sky130_fd_sc_hd__a22o_1 _16653_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_06017_),
    .B2(_05185_),
    .X(_06041_));
 sky130_fd_sc_hd__a21oi_1 _16654_ (.A1(_06018_),
    .A2(_06033_),
    .B1(net267),
    .Y(_06042_));
 sky130_fd_sc_hd__o21ai_4 _16655_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_06036_),
    .Y(_06043_));
 sky130_fd_sc_hd__o21ai_4 _16656_ (.A1(_06041_),
    .A2(_06034_),
    .B1(_06040_),
    .Y(_06044_));
 sky130_fd_sc_hd__o211ai_4 _16657_ (.A1(_05527_),
    .A2(_05539_),
    .B1(_05792_),
    .C1(_05531_),
    .Y(_06045_));
 sky130_fd_sc_hd__o22ai_2 _16658_ (.A1(_05790_),
    .A2(_05782_),
    .B1(_05788_),
    .B2(_05794_),
    .Y(_06046_));
 sky130_fd_sc_hd__o21ai_2 _16659_ (.A1(net293),
    .A2(_05784_),
    .B1(_06045_),
    .Y(_06047_));
 sky130_fd_sc_hd__o2111ai_4 _16660_ (.A1(net293),
    .A2(_05784_),
    .B1(_06040_),
    .C1(_06043_),
    .D1(_06045_),
    .Y(_06049_));
 sky130_fd_sc_hd__o311a_1 _16661_ (.A1(net295),
    .A2(_05782_),
    .A3(_05783_),
    .B1(_05797_),
    .C1(_06044_),
    .X(_06050_));
 sky130_fd_sc_hd__o211ai_2 _16662_ (.A1(_05794_),
    .A2(_05793_),
    .B1(_05792_),
    .C1(_06044_),
    .Y(_06051_));
 sky130_fd_sc_hd__o22ai_2 _16663_ (.A1(net402),
    .A2(net400),
    .B1(_06044_),
    .B2(_06047_),
    .Y(_06052_));
 sky130_fd_sc_hd__o211ai_2 _16664_ (.A1(net402),
    .A2(net400),
    .B1(_06049_),
    .C1(_06051_),
    .Y(_06053_));
 sky130_fd_sc_hd__o22ai_4 _16665_ (.A1(net388),
    .A2(_06035_),
    .B1(_06052_),
    .B2(_06050_),
    .Y(_06054_));
 sky130_fd_sc_hd__a2bb2oi_2 _16666_ (.A1_N(_05242_),
    .A2_N(net317),
    .B1(_06039_),
    .B2(_06053_),
    .Y(_06055_));
 sky130_fd_sc_hd__o21ai_2 _16667_ (.A1(_05242_),
    .A2(net317),
    .B1(_06054_),
    .Y(_06056_));
 sky130_fd_sc_hd__a31oi_2 _16668_ (.A1(net388),
    .A2(_06049_),
    .A3(_06051_),
    .B1(net293),
    .Y(_06057_));
 sky130_fd_sc_hd__a31o_1 _16669_ (.A1(net388),
    .A2(_06049_),
    .A3(_06051_),
    .B1(net293),
    .X(_06058_));
 sky130_fd_sc_hd__and3_2 _16670_ (.A(_06053_),
    .B(net295),
    .C(_06039_),
    .X(_06060_));
 sky130_fd_sc_hd__o211ai_1 _16671_ (.A1(net388),
    .A2(_06035_),
    .B1(net295),
    .C1(_06053_),
    .Y(_06061_));
 sky130_fd_sc_hd__a21oi_1 _16672_ (.A1(_06039_),
    .A2(_06057_),
    .B1(_06055_),
    .Y(_06062_));
 sky130_fd_sc_hd__a21oi_1 _16673_ (.A1(_05804_),
    .A2(_05806_),
    .B1(_05801_),
    .Y(_06063_));
 sky130_fd_sc_hd__o21ai_2 _16674_ (.A1(_05803_),
    .A2(_05805_),
    .B1(_05802_),
    .Y(_06064_));
 sky130_fd_sc_hd__a21oi_1 _16675_ (.A1(_06056_),
    .A2(_06061_),
    .B1(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__o21ai_1 _16676_ (.A1(_06055_),
    .A2(_06060_),
    .B1(_06063_),
    .Y(_06066_));
 sky130_fd_sc_hd__o211a_1 _16677_ (.A1(_06058_),
    .A2(_06038_),
    .B1(_06056_),
    .C1(_06064_),
    .X(_06067_));
 sky130_fd_sc_hd__o211ai_2 _16678_ (.A1(_06058_),
    .A2(_06038_),
    .B1(_06056_),
    .C1(_06064_),
    .Y(_06068_));
 sky130_fd_sc_hd__o22ai_2 _16679_ (.A1(net384),
    .A2(net383),
    .B1(_06065_),
    .B2(_06067_),
    .Y(_06069_));
 sky130_fd_sc_hd__and3_1 _16680_ (.A(_05687_),
    .B(_05709_),
    .C(_06054_),
    .X(_06071_));
 sky130_fd_sc_hd__a211o_1 _16681_ (.A1(_06039_),
    .A2(_06053_),
    .B1(net384),
    .C1(net383),
    .X(_06072_));
 sky130_fd_sc_hd__nand3_1 _16682_ (.A(_06066_),
    .B(_06068_),
    .C(net359),
    .Y(_06073_));
 sky130_fd_sc_hd__o31a_2 _16683_ (.A1(_05731_),
    .A2(_06065_),
    .A3(_06067_),
    .B1(_06072_),
    .X(_06074_));
 sky130_fd_sc_hd__o311a_1 _16684_ (.A1(net384),
    .A2(_06054_),
    .A3(net383),
    .B1(_06848_),
    .C1(_06069_),
    .X(_06075_));
 sky130_fd_sc_hd__or3_2 _16685_ (.A(net379),
    .B(net378),
    .C(_06074_),
    .X(_06076_));
 sky130_fd_sc_hd__a2bb2oi_1 _16686_ (.A1_N(net339),
    .A2_N(_04184_),
    .B1(_06072_),
    .B2(_06073_),
    .Y(_06077_));
 sky130_fd_sc_hd__o221ai_4 _16687_ (.A1(net339),
    .A2(_04184_),
    .B1(_06054_),
    .B2(net359),
    .C1(_06069_),
    .Y(_06078_));
 sky130_fd_sc_hd__a31oi_1 _16688_ (.A1(_06066_),
    .A2(_06068_),
    .A3(net359),
    .B1(net298),
    .Y(_06079_));
 sky130_fd_sc_hd__a31o_1 _16689_ (.A1(_06066_),
    .A2(_06068_),
    .A3(net359),
    .B1(net298),
    .X(_06080_));
 sky130_fd_sc_hd__o311a_1 _16690_ (.A1(_05731_),
    .A2(_06065_),
    .A3(_06067_),
    .B1(_06072_),
    .C1(net299),
    .X(_06082_));
 sky130_fd_sc_hd__a21oi_2 _16691_ (.A1(_06072_),
    .A2(_06079_),
    .B1(_06077_),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_4 _16692_ (.A1(_06071_),
    .A2(_06080_),
    .B1(_06078_),
    .Y(_06084_));
 sky130_fd_sc_hd__a22oi_4 _16693_ (.A1(_02148_),
    .A2(_05811_),
    .B1(_05828_),
    .B2(_05826_),
    .Y(_06085_));
 sky130_fd_sc_hd__o2bb2ai_2 _16694_ (.A1_N(_02148_),
    .A2_N(_05811_),
    .B1(_05830_),
    .B2(_05825_),
    .Y(_06086_));
 sky130_fd_sc_hd__a21oi_4 _16695_ (.A1(_05813_),
    .A2(_05833_),
    .B1(_06084_),
    .Y(_06087_));
 sky130_fd_sc_hd__nand2_2 _16696_ (.A(_06083_),
    .B(_06086_),
    .Y(_06088_));
 sky130_fd_sc_hd__o21ai_1 _16697_ (.A1(_06077_),
    .A2(_06082_),
    .B1(_06085_),
    .Y(_06089_));
 sky130_fd_sc_hd__o22ai_4 _16698_ (.A1(net379),
    .A2(net378),
    .B1(_06086_),
    .B2(_06083_),
    .Y(_06090_));
 sky130_fd_sc_hd__nand3_1 _16699_ (.A(_06088_),
    .B(_06089_),
    .C(net357),
    .Y(_06091_));
 sky130_fd_sc_hd__o22a_1 _16700_ (.A1(net357),
    .A2(_06074_),
    .B1(_06087_),
    .B2(_06090_),
    .X(_06093_));
 sky130_fd_sc_hd__o21ai_4 _16701_ (.A1(_06087_),
    .A2(_06090_),
    .B1(_06076_),
    .Y(_06094_));
 sky130_fd_sc_hd__a2bb2oi_2 _16702_ (.A1_N(_02049_),
    .A2_N(net342),
    .B1(_06076_),
    .B2(_06091_),
    .Y(_06095_));
 sky130_fd_sc_hd__o21ai_4 _16703_ (.A1(_02049_),
    .A2(net342),
    .B1(_06094_),
    .Y(_06096_));
 sky130_fd_sc_hd__a31o_1 _16704_ (.A1(_06088_),
    .A2(_06089_),
    .A3(net357),
    .B1(_02148_),
    .X(_06097_));
 sky130_fd_sc_hd__o221a_2 _16705_ (.A1(net357),
    .A2(_06074_),
    .B1(_06087_),
    .B2(_06090_),
    .C1(_02137_),
    .X(_06098_));
 sky130_fd_sc_hd__o221ai_4 _16706_ (.A1(net357),
    .A2(_06074_),
    .B1(_06087_),
    .B2(_06090_),
    .C1(_02137_),
    .Y(_06099_));
 sky130_fd_sc_hd__o21ai_2 _16707_ (.A1(net320),
    .A2(_05839_),
    .B1(_05849_),
    .Y(_06100_));
 sky130_fd_sc_hd__o22a_1 _16708_ (.A1(_05843_),
    .A2(_05837_),
    .B1(_05848_),
    .B2(_05846_),
    .X(_06101_));
 sky130_fd_sc_hd__o22ai_4 _16709_ (.A1(_05843_),
    .A2(_05837_),
    .B1(_05848_),
    .B2(_05846_),
    .Y(_06102_));
 sky130_fd_sc_hd__o211ai_1 _16710_ (.A1(_06075_),
    .A2(_06097_),
    .B1(_06102_),
    .C1(_06096_),
    .Y(_06104_));
 sky130_fd_sc_hd__o21ai_1 _16711_ (.A1(_06095_),
    .A2(_06098_),
    .B1(_06101_),
    .Y(_06105_));
 sky130_fd_sc_hd__o211ai_4 _16712_ (.A1(_06075_),
    .A2(_06097_),
    .B1(_06096_),
    .C1(_06101_),
    .Y(_06106_));
 sky130_fd_sc_hd__o21ai_2 _16713_ (.A1(_06095_),
    .A2(_06098_),
    .B1(_06102_),
    .Y(_06107_));
 sky130_fd_sc_hd__nand3_2 _16714_ (.A(_06105_),
    .B(net356),
    .C(_06104_),
    .Y(_06108_));
 sky130_fd_sc_hd__a21oi_1 _16715_ (.A1(_06076_),
    .A2(_06091_),
    .B1(net356),
    .Y(_06109_));
 sky130_fd_sc_hd__or3_1 _16716_ (.A(net372),
    .B(net371),
    .C(_06093_),
    .X(_06110_));
 sky130_fd_sc_hd__o211ai_4 _16717_ (.A1(net372),
    .A2(net371),
    .B1(_06106_),
    .C1(_06107_),
    .Y(_06111_));
 sky130_fd_sc_hd__o31a_1 _16718_ (.A1(net372),
    .A2(net371),
    .A3(_06093_),
    .B1(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__o211a_2 _16719_ (.A1(_06094_),
    .A2(net356),
    .B1(_08732_),
    .C1(_06108_),
    .X(_06113_));
 sky130_fd_sc_hd__a211o_1 _16720_ (.A1(_06110_),
    .A2(_06111_),
    .B1(net353),
    .C1(net352),
    .X(_06115_));
 sky130_fd_sc_hd__a311oi_4 _16721_ (.A1(_06106_),
    .A2(_06107_),
    .A3(net356),
    .B1(_06109_),
    .C1(net319),
    .Y(_06116_));
 sky130_fd_sc_hd__nand3_4 _16722_ (.A(_06111_),
    .B(net320),
    .C(_06110_),
    .Y(_06117_));
 sky130_fd_sc_hd__o211a_1 _16723_ (.A1(_06094_),
    .A2(net356),
    .B1(net319),
    .C1(_06108_),
    .X(_06118_));
 sky130_fd_sc_hd__o211ai_4 _16724_ (.A1(_06094_),
    .A2(net356),
    .B1(net319),
    .C1(_06108_),
    .Y(_06119_));
 sky130_fd_sc_hd__o21a_1 _16725_ (.A1(_12888_),
    .A2(_05854_),
    .B1(_05859_),
    .X(_06120_));
 sky130_fd_sc_hd__a31oi_2 _16726_ (.A1(_05842_),
    .A2(_05853_),
    .A3(_12888_),
    .B1(_05859_),
    .Y(_06121_));
 sky130_fd_sc_hd__o21ai_1 _16727_ (.A1(_05859_),
    .A2(_05861_),
    .B1(_05865_),
    .Y(_06122_));
 sky130_fd_sc_hd__a21oi_1 _16728_ (.A1(_05863_),
    .A2(_05858_),
    .B1(_05864_),
    .Y(_06123_));
 sky130_fd_sc_hd__a21oi_2 _16729_ (.A1(_06117_),
    .A2(_06119_),
    .B1(_06122_),
    .Y(_06124_));
 sky130_fd_sc_hd__o2bb2ai_4 _16730_ (.A1_N(_06117_),
    .A2_N(_06119_),
    .B1(_06120_),
    .B2(_05861_),
    .Y(_06126_));
 sky130_fd_sc_hd__o211ai_4 _16731_ (.A1(_05864_),
    .A2(_06121_),
    .B1(_06119_),
    .C1(_06117_),
    .Y(_06127_));
 sky130_fd_sc_hd__o21ai_2 _16732_ (.A1(net353),
    .A2(net352),
    .B1(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__nand3_1 _16733_ (.A(_06126_),
    .B(_06127_),
    .C(_08721_),
    .Y(_06129_));
 sky130_fd_sc_hd__a31oi_4 _16734_ (.A1(_06126_),
    .A2(_06127_),
    .A3(_08721_),
    .B1(_06113_),
    .Y(_06130_));
 sky130_fd_sc_hd__o22ai_4 _16735_ (.A1(_08721_),
    .A2(_06112_),
    .B1(_06124_),
    .B2(_06128_),
    .Y(_06131_));
 sky130_fd_sc_hd__o221a_1 _16736_ (.A1(_08721_),
    .A2(_06112_),
    .B1(_06124_),
    .B2(_06128_),
    .C1(_09840_),
    .X(_06132_));
 sky130_fd_sc_hd__o21ai_1 _16737_ (.A1(_05620_),
    .A2(_05878_),
    .B1(_05877_),
    .Y(_06133_));
 sky130_fd_sc_hd__a31oi_1 _16738_ (.A1(net331),
    .A2(_05871_),
    .A3(_05872_),
    .B1(_05880_),
    .Y(_06134_));
 sky130_fd_sc_hd__a21oi_2 _16739_ (.A1(_05875_),
    .A2(_05879_),
    .B1(_05876_),
    .Y(_06135_));
 sky130_fd_sc_hd__a311oi_4 _16740_ (.A1(_06126_),
    .A2(_06127_),
    .A3(_08721_),
    .B1(net325),
    .C1(_06113_),
    .Y(_06137_));
 sky130_fd_sc_hd__a311o_1 _16741_ (.A1(_06126_),
    .A2(_06127_),
    .A3(_08721_),
    .B1(net325),
    .C1(_06113_),
    .X(_06138_));
 sky130_fd_sc_hd__a2bb2oi_1 _16742_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_06115_),
    .B2(_06129_),
    .Y(_06139_));
 sky130_fd_sc_hd__o21ai_1 _16743_ (.A1(_12845_),
    .A2(_12856_),
    .B1(_06131_),
    .Y(_06140_));
 sky130_fd_sc_hd__nand3_1 _16744_ (.A(_06135_),
    .B(_06138_),
    .C(_06140_),
    .Y(_06141_));
 sky130_fd_sc_hd__o22ai_2 _16745_ (.A1(_05876_),
    .A2(_06134_),
    .B1(_06137_),
    .B2(_06139_),
    .Y(_06142_));
 sky130_fd_sc_hd__nand3_1 _16746_ (.A(_06141_),
    .B(_06142_),
    .C(net337),
    .Y(_06143_));
 sky130_fd_sc_hd__or3_2 _16747_ (.A(net350),
    .B(net349),
    .C(_06130_),
    .X(_06144_));
 sky130_fd_sc_hd__o221ai_4 _16748_ (.A1(_05874_),
    .A2(net330),
    .B1(_12888_),
    .B2(_06130_),
    .C1(_06133_),
    .Y(_06145_));
 sky130_fd_sc_hd__o21ai_1 _16749_ (.A1(_06137_),
    .A2(_06139_),
    .B1(_06135_),
    .Y(_06146_));
 sky130_fd_sc_hd__o221ai_4 _16750_ (.A1(net350),
    .A2(net349),
    .B1(_06137_),
    .B2(_06145_),
    .C1(_06146_),
    .Y(_06148_));
 sky130_fd_sc_hd__a31o_1 _16751_ (.A1(_06141_),
    .A2(_06142_),
    .A3(net337),
    .B1(_06132_),
    .X(_06149_));
 sky130_fd_sc_hd__nand2_1 _16752_ (.A(_11079_),
    .B(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__o211ai_4 _16753_ (.A1(_06131_),
    .A2(net337),
    .B1(net330),
    .C1(_06143_),
    .Y(_06151_));
 sky130_fd_sc_hd__and3_1 _16754_ (.A(_06148_),
    .B(net331),
    .C(_06144_),
    .X(_06152_));
 sky130_fd_sc_hd__nand3_4 _16755_ (.A(_06148_),
    .B(net331),
    .C(_06144_),
    .Y(_06153_));
 sky130_fd_sc_hd__o21a_1 _16756_ (.A1(_10015_),
    .A2(_05887_),
    .B1(_05890_),
    .X(_06154_));
 sky130_fd_sc_hd__o32a_1 _16757_ (.A1(_09971_),
    .A2(net363),
    .A3(_05887_),
    .B1(_05890_),
    .B2(_05892_),
    .X(_06155_));
 sky130_fd_sc_hd__o32ai_2 _16758_ (.A1(_09971_),
    .A2(net363),
    .A3(_05887_),
    .B1(_05890_),
    .B2(_05892_),
    .Y(_06156_));
 sky130_fd_sc_hd__a21oi_1 _16759_ (.A1(_06151_),
    .A2(_06153_),
    .B1(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__o2bb2ai_2 _16760_ (.A1_N(_06151_),
    .A2_N(_06153_),
    .B1(_06154_),
    .B2(_05892_),
    .Y(_06159_));
 sky130_fd_sc_hd__o2111a_1 _16761_ (.A1(_05888_),
    .A2(_05891_),
    .B1(_05893_),
    .C1(_06151_),
    .D1(_06153_),
    .X(_06160_));
 sky130_fd_sc_hd__o2111ai_4 _16762_ (.A1(_05888_),
    .A2(_05891_),
    .B1(_05893_),
    .C1(_06151_),
    .D1(_06153_),
    .Y(_06161_));
 sky130_fd_sc_hd__o22ai_2 _16763_ (.A1(net347),
    .A2(net346),
    .B1(_06157_),
    .B2(_06160_),
    .Y(_06162_));
 sky130_fd_sc_hd__o211a_2 _16764_ (.A1(_06131_),
    .A2(net337),
    .B1(_11079_),
    .C1(_06143_),
    .X(_06163_));
 sky130_fd_sc_hd__a311o_1 _16765_ (.A1(_06141_),
    .A2(_06142_),
    .A3(net337),
    .B1(net334),
    .C1(_06132_),
    .X(_06164_));
 sky130_fd_sc_hd__nand3_2 _16766_ (.A(_06159_),
    .B(_06161_),
    .C(net334),
    .Y(_06165_));
 sky130_fd_sc_hd__a31o_1 _16767_ (.A1(_06159_),
    .A2(_06161_),
    .A3(net334),
    .B1(_06163_),
    .X(_06166_));
 sky130_fd_sc_hd__a311o_1 _16768_ (.A1(_06159_),
    .A2(_06161_),
    .A3(net334),
    .B1(_06163_),
    .C1(net313),
    .X(_06167_));
 sky130_fd_sc_hd__a2bb2oi_4 _16769_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_06164_),
    .B2(_06165_),
    .Y(_06168_));
 sky130_fd_sc_hd__o211ai_4 _16770_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_06150_),
    .C1(_06162_),
    .Y(_06170_));
 sky130_fd_sc_hd__a31o_1 _16771_ (.A1(_06159_),
    .A2(_06161_),
    .A3(net334),
    .B1(net348),
    .X(_06171_));
 sky130_fd_sc_hd__o221a_1 _16772_ (.A1(_09971_),
    .A2(net363),
    .B1(net334),
    .B2(_06149_),
    .C1(_06165_),
    .X(_06172_));
 sky130_fd_sc_hd__a32oi_4 _16773_ (.A1(_05897_),
    .A2(_05899_),
    .A3(_08907_),
    .B1(_05656_),
    .B2(_05657_),
    .Y(_06173_));
 sky130_fd_sc_hd__a21oi_2 _16774_ (.A1(_05910_),
    .A2(_05902_),
    .B1(_05911_),
    .Y(_06174_));
 sky130_fd_sc_hd__a21o_1 _16775_ (.A1(_05910_),
    .A2(_05902_),
    .B1(_05911_),
    .X(_06175_));
 sky130_fd_sc_hd__o21ai_2 _16776_ (.A1(_06168_),
    .A2(_06172_),
    .B1(_06174_),
    .Y(_06176_));
 sky130_fd_sc_hd__o22a_1 _16777_ (.A1(net348),
    .A2(_06166_),
    .B1(_06173_),
    .B2(_05911_),
    .X(_06177_));
 sky130_fd_sc_hd__o22ai_2 _16778_ (.A1(net348),
    .A2(_06166_),
    .B1(_06173_),
    .B2(_05911_),
    .Y(_06178_));
 sky130_fd_sc_hd__o221ai_4 _16779_ (.A1(_05911_),
    .A2(_06173_),
    .B1(_06163_),
    .B2(_06171_),
    .C1(_06170_),
    .Y(_06179_));
 sky130_fd_sc_hd__o211ai_1 _16780_ (.A1(_06163_),
    .A2(_06171_),
    .B1(_06170_),
    .C1(_06174_),
    .Y(_06181_));
 sky130_fd_sc_hd__o21ai_1 _16781_ (.A1(_06168_),
    .A2(_06172_),
    .B1(_06175_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand3_2 _16782_ (.A(_06182_),
    .B(net313),
    .C(_06181_),
    .Y(_06183_));
 sky130_fd_sc_hd__and3_1 _16783_ (.A(_12703_),
    .B(_06150_),
    .C(_06162_),
    .X(_06184_));
 sky130_fd_sc_hd__a211o_2 _16784_ (.A1(_06164_),
    .A2(_06165_),
    .B1(net328),
    .C1(_12681_),
    .X(_06185_));
 sky130_fd_sc_hd__nand3_2 _16785_ (.A(_06176_),
    .B(_06179_),
    .C(net313),
    .Y(_06186_));
 sky130_fd_sc_hd__a311oi_4 _16786_ (.A1(_06176_),
    .A2(_06179_),
    .A3(net313),
    .B1(_06184_),
    .C1(_08918_),
    .Y(_06187_));
 sky130_fd_sc_hd__o211ai_2 _16787_ (.A1(_08863_),
    .A2(net366),
    .B1(_06185_),
    .C1(_06186_),
    .Y(_06188_));
 sky130_fd_sc_hd__a2bb2oi_4 _16788_ (.A1_N(_08819_),
    .A2_N(net367),
    .B1(_06185_),
    .B2(_06186_),
    .Y(_06189_));
 sky130_fd_sc_hd__o211ai_4 _16789_ (.A1(_08819_),
    .A2(net367),
    .B1(_06167_),
    .C1(_06183_),
    .Y(_06190_));
 sky130_fd_sc_hd__nand3_4 _16790_ (.A(_06006_),
    .B(_06188_),
    .C(_06190_),
    .Y(_06192_));
 sky130_fd_sc_hd__o22ai_4 _16791_ (.A1(_05918_),
    .A2(_06005_),
    .B1(_06187_),
    .B2(_06189_),
    .Y(_06193_));
 sky130_fd_sc_hd__nand3_2 _16792_ (.A(_06193_),
    .B(net310),
    .C(_06192_),
    .Y(_06194_));
 sky130_fd_sc_hd__o311a_2 _16793_ (.A1(net328),
    .A2(_12681_),
    .A3(_06166_),
    .B1(_06183_),
    .C1(_00066_),
    .X(_06195_));
 sky130_fd_sc_hd__a211o_2 _16794_ (.A1(_06185_),
    .A2(_06186_),
    .B1(net324),
    .C1(net322),
    .X(_06196_));
 sky130_fd_sc_hd__a31o_4 _16795_ (.A1(_06193_),
    .A2(net310),
    .A3(_06192_),
    .B1(_06195_),
    .X(_06197_));
 sky130_fd_sc_hd__o221a_1 _16796_ (.A1(_05680_),
    .A2(_06332_),
    .B1(_07033_),
    .B2(_05926_),
    .C1(_05693_),
    .X(_06198_));
 sky130_fd_sc_hd__a21oi_2 _16797_ (.A1(_05684_),
    .A2(_05693_),
    .B1(_05930_),
    .Y(_06199_));
 sky130_fd_sc_hd__o21ai_2 _16798_ (.A1(_05929_),
    .A2(_05930_),
    .B1(_05933_),
    .Y(_06200_));
 sky130_fd_sc_hd__a311oi_4 _16799_ (.A1(_06193_),
    .A2(net310),
    .A3(_06192_),
    .B1(_06195_),
    .C1(_07899_),
    .Y(_06201_));
 sky130_fd_sc_hd__o211ai_2 _16800_ (.A1(net369),
    .A2(_07866_),
    .B1(_06194_),
    .C1(_06196_),
    .Y(_06202_));
 sky130_fd_sc_hd__a22oi_4 _16801_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_06194_),
    .B2(_06196_),
    .Y(_06203_));
 sky130_fd_sc_hd__a22o_1 _16802_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_06194_),
    .B2(_06196_),
    .X(_06204_));
 sky130_fd_sc_hd__o211ai_1 _16803_ (.A1(_05930_),
    .A2(_06198_),
    .B1(_06202_),
    .C1(_06204_),
    .Y(_06205_));
 sky130_fd_sc_hd__o22ai_1 _16804_ (.A1(_05932_),
    .A2(_06199_),
    .B1(_06201_),
    .B2(_06203_),
    .Y(_06206_));
 sky130_fd_sc_hd__nand3_2 _16805_ (.A(_06205_),
    .B(_06206_),
    .C(_01962_),
    .Y(_06207_));
 sky130_fd_sc_hd__a211o_2 _16806_ (.A1(_06194_),
    .A2(_06196_),
    .B1(net306),
    .C1(net303),
    .X(_06208_));
 sky130_fd_sc_hd__o22a_1 _16807_ (.A1(_07899_),
    .A2(_06197_),
    .B1(_06199_),
    .B2(_05932_),
    .X(_06209_));
 sky130_fd_sc_hd__o221ai_2 _16808_ (.A1(_07899_),
    .A2(_06197_),
    .B1(_06199_),
    .B2(_05932_),
    .C1(_06204_),
    .Y(_06210_));
 sky130_fd_sc_hd__o22ai_1 _16809_ (.A1(_05930_),
    .A2(_06198_),
    .B1(_06201_),
    .B2(_06203_),
    .Y(_06211_));
 sky130_fd_sc_hd__nand3_2 _16810_ (.A(_06210_),
    .B(_06211_),
    .C(_01962_),
    .Y(_06213_));
 sky130_fd_sc_hd__o21a_2 _16811_ (.A1(net280),
    .A2(_06197_),
    .B1(_06207_),
    .X(_06214_));
 sky130_fd_sc_hd__a21oi_2 _16812_ (.A1(_05943_),
    .A2(_05947_),
    .B1(_05944_),
    .Y(_06215_));
 sky130_fd_sc_hd__o32ai_4 _16813_ (.A1(_06332_),
    .A2(_05927_),
    .A3(_05937_),
    .B1(_05942_),
    .B2(_05946_),
    .Y(_06216_));
 sky130_fd_sc_hd__and3_1 _16814_ (.A(_06213_),
    .B(_07033_),
    .C(_06208_),
    .X(_06217_));
 sky130_fd_sc_hd__o211ai_4 _16815_ (.A1(_06989_),
    .A2(_07011_),
    .B1(_06208_),
    .C1(_06213_),
    .Y(_06218_));
 sky130_fd_sc_hd__o211a_1 _16816_ (.A1(_06197_),
    .A2(net280),
    .B1(_07044_),
    .C1(_06207_),
    .X(_06219_));
 sky130_fd_sc_hd__o211ai_4 _16817_ (.A1(_06197_),
    .A2(net280),
    .B1(_07044_),
    .C1(_06207_),
    .Y(_06220_));
 sky130_fd_sc_hd__a21oi_4 _16818_ (.A1(_06218_),
    .A2(_06220_),
    .B1(_06215_),
    .Y(_06221_));
 sky130_fd_sc_hd__a31o_2 _16819_ (.A1(_06215_),
    .A2(_06218_),
    .A3(_06220_),
    .B1(_04040_),
    .X(_06222_));
 sky130_fd_sc_hd__nand3_1 _16820_ (.A(_06216_),
    .B(_06218_),
    .C(_06220_),
    .Y(_06224_));
 sky130_fd_sc_hd__a21o_1 _16821_ (.A1(_06218_),
    .A2(_06220_),
    .B1(_06216_),
    .X(_06225_));
 sky130_fd_sc_hd__nand3_1 _16822_ (.A(_06225_),
    .B(net275),
    .C(_06224_),
    .Y(_06226_));
 sky130_fd_sc_hd__a211o_1 _16823_ (.A1(_06208_),
    .A2(_06213_),
    .B1(net301),
    .C1(net300),
    .X(_06227_));
 sky130_fd_sc_hd__o22ai_4 _16824_ (.A1(net275),
    .A2(_06214_),
    .B1(_06221_),
    .B2(_06222_),
    .Y(_06228_));
 sky130_fd_sc_hd__o221a_1 _16825_ (.A1(net275),
    .A2(_06214_),
    .B1(_06221_),
    .B2(_06222_),
    .C1(_06343_),
    .X(_06229_));
 sky130_fd_sc_hd__o221ai_4 _16826_ (.A1(net275),
    .A2(_06214_),
    .B1(_06221_),
    .B2(_06222_),
    .C1(_06343_),
    .Y(_06230_));
 sky130_fd_sc_hd__nand3_2 _16827_ (.A(_06226_),
    .B(_06227_),
    .C(_06332_),
    .Y(_06231_));
 sky130_fd_sc_hd__o21ai_1 _16828_ (.A1(_05941_),
    .A2(_05953_),
    .B1(_05960_),
    .Y(_06232_));
 sky130_fd_sc_hd__a22oi_1 _16829_ (.A1(_05955_),
    .A2(_05956_),
    .B1(_05959_),
    .B2(_05862_),
    .Y(_06233_));
 sky130_fd_sc_hd__o2bb2ai_2 _16830_ (.A1_N(_06230_),
    .A2_N(_06231_),
    .B1(_06233_),
    .B2(_05962_),
    .Y(_06235_));
 sky130_fd_sc_hd__a22oi_2 _16831_ (.A1(_06228_),
    .A2(_06332_),
    .B1(_05964_),
    .B2(_06232_),
    .Y(_06236_));
 sky130_fd_sc_hd__o211ai_1 _16832_ (.A1(_05963_),
    .A2(_05957_),
    .B1(_05960_),
    .C1(_06231_),
    .Y(_06237_));
 sky130_fd_sc_hd__o2111ai_4 _16833_ (.A1(_05963_),
    .A2(_05957_),
    .B1(_05960_),
    .C1(_06230_),
    .D1(_06231_),
    .Y(_06238_));
 sky130_fd_sc_hd__nand3_1 _16834_ (.A(_06235_),
    .B(_06238_),
    .C(net274),
    .Y(_06239_));
 sky130_fd_sc_hd__o221a_2 _16835_ (.A1(net275),
    .A2(_06214_),
    .B1(_06221_),
    .B2(_06222_),
    .C1(_05234_),
    .X(_06240_));
 sky130_fd_sc_hd__or3_1 _16836_ (.A(net297),
    .B(_05232_),
    .C(_06228_),
    .X(_06241_));
 sky130_fd_sc_hd__a31o_1 _16837_ (.A1(_06235_),
    .A2(_06238_),
    .A3(net274),
    .B1(_06240_),
    .X(_06242_));
 sky130_fd_sc_hd__a31oi_2 _16838_ (.A1(_06235_),
    .A2(_06238_),
    .A3(net274),
    .B1(_06240_),
    .Y(_06243_));
 sky130_fd_sc_hd__nand4_4 _16839_ (.A(_05739_),
    .B(_05741_),
    .C(_05966_),
    .D(_05968_),
    .Y(_06244_));
 sky130_fd_sc_hd__o211ai_4 _16840_ (.A1(net387),
    .A2(_05970_),
    .B1(_05978_),
    .C1(_06244_),
    .Y(_06246_));
 sky130_fd_sc_hd__o2111ai_4 _16841_ (.A1(net387),
    .A2(_05970_),
    .B1(_05978_),
    .C1(_05851_),
    .D1(_06244_),
    .Y(_06247_));
 sky130_fd_sc_hd__o21ai_1 _16842_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_06246_),
    .Y(_06248_));
 sky130_fd_sc_hd__and4_1 _16843_ (.A(_06248_),
    .B(_06242_),
    .C(_05485_),
    .D(_06247_),
    .X(_06249_));
 sky130_fd_sc_hd__nand4_1 _16844_ (.A(_06248_),
    .B(_06242_),
    .C(_05485_),
    .D(_06247_),
    .Y(_06250_));
 sky130_fd_sc_hd__a31oi_1 _16845_ (.A1(_06248_),
    .A2(_05485_),
    .A3(_06247_),
    .B1(_06242_),
    .Y(_06251_));
 sky130_fd_sc_hd__a31o_1 _16846_ (.A1(_06248_),
    .A2(_05485_),
    .A3(_06247_),
    .B1(_06242_),
    .X(_06252_));
 sky130_fd_sc_hd__and3_2 _16847_ (.A(_06242_),
    .B(_05484_),
    .C(_05482_),
    .X(_06253_));
 sky130_fd_sc_hd__a22oi_1 _16848_ (.A1(_05774_),
    .A2(_05796_),
    .B1(_06239_),
    .B2(_06241_),
    .Y(_06254_));
 sky130_fd_sc_hd__a31oi_1 _16849_ (.A1(_06235_),
    .A2(_06238_),
    .A3(net274),
    .B1(_05862_),
    .Y(_06255_));
 sky130_fd_sc_hd__a31o_1 _16850_ (.A1(_06235_),
    .A2(_06238_),
    .A3(net274),
    .B1(_05862_),
    .X(_06257_));
 sky130_fd_sc_hd__o311a_1 _16851_ (.A1(net297),
    .A2(_05232_),
    .A3(_06228_),
    .B1(_05851_),
    .C1(_06239_),
    .X(_06258_));
 sky130_fd_sc_hd__o221ai_4 _16852_ (.A1(_05851_),
    .A2(_06243_),
    .B1(_06240_),
    .B2(_06257_),
    .C1(_06246_),
    .Y(_06259_));
 sky130_fd_sc_hd__a22oi_1 _16853_ (.A1(_06255_),
    .A2(_06241_),
    .B1(_06242_),
    .B2(_05862_),
    .Y(_06260_));
 sky130_fd_sc_hd__o21bai_1 _16854_ (.A1(_06254_),
    .A2(_06258_),
    .B1_N(_06246_),
    .Y(_06261_));
 sky130_fd_sc_hd__o221a_2 _16855_ (.A1(_05481_),
    .A2(net269),
    .B1(_06246_),
    .B2(_06260_),
    .C1(_06259_),
    .X(_06262_));
 sky130_fd_sc_hd__a31oi_4 _16856_ (.A1(_06261_),
    .A2(_05485_),
    .A3(_06259_),
    .B1(_06253_),
    .Y(_06263_));
 sky130_fd_sc_hd__o211ai_4 _16857_ (.A1(net398),
    .A2(net397),
    .B1(_05982_),
    .C1(_05986_),
    .Y(_06264_));
 sky130_fd_sc_hd__o22ai_4 _16858_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_05981_),
    .B2(_05985_),
    .Y(_06265_));
 sky130_fd_sc_hd__nand3_1 _16859_ (.A(_06265_),
    .B(net241),
    .C(_06264_),
    .Y(_06266_));
 sky130_fd_sc_hd__a31o_1 _16860_ (.A1(_06265_),
    .A2(net241),
    .A3(_06264_),
    .B1(_06263_),
    .X(_06268_));
 sky130_fd_sc_hd__nand4_2 _16861_ (.A(_06263_),
    .B(_06264_),
    .C(_06265_),
    .D(net241),
    .Y(_06269_));
 sky130_fd_sc_hd__o2111ai_4 _16862_ (.A1(_06253_),
    .A2(_06262_),
    .B1(net241),
    .C1(_06264_),
    .D1(_06265_),
    .Y(_06270_));
 sky130_fd_sc_hd__o21ai_2 _16863_ (.A1(_06249_),
    .A2(_06251_),
    .B1(_06266_),
    .Y(_06271_));
 sky130_fd_sc_hd__nand2_1 _16864_ (.A(_06270_),
    .B(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__and3_1 _16865_ (.A(_06271_),
    .B(net403),
    .C(_06270_),
    .X(_06273_));
 sky130_fd_sc_hd__nand3_2 _16866_ (.A(_06271_),
    .B(net403),
    .C(_06270_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand3_4 _16867_ (.A(_05250_),
    .B(_06268_),
    .C(_06269_),
    .Y(_06275_));
 sky130_fd_sc_hd__a21oi_1 _16868_ (.A1(_06274_),
    .A2(_06275_),
    .B1(_05999_),
    .Y(_06276_));
 sky130_fd_sc_hd__o21ai_2 _16869_ (.A1(_03289_),
    .A2(_05988_),
    .B1(_06274_),
    .Y(_06277_));
 sky130_fd_sc_hd__o211a_1 _16870_ (.A1(_03289_),
    .A2(_05988_),
    .B1(_06274_),
    .C1(_06275_),
    .X(_06279_));
 sky130_fd_sc_hd__o2bb2ai_1 _16871_ (.A1_N(_06274_),
    .A2_N(_06275_),
    .B1(_03289_),
    .B2(_05988_),
    .Y(_06280_));
 sky130_fd_sc_hd__a31o_1 _16872_ (.A1(_05250_),
    .A2(_06268_),
    .A3(_06269_),
    .B1(_05999_),
    .X(_06281_));
 sky130_fd_sc_hd__o211ai_4 _16873_ (.A1(_06273_),
    .A2(_06281_),
    .B1(_06280_),
    .C1(_05996_),
    .Y(_06282_));
 sky130_fd_sc_hd__or3_2 _16874_ (.A(net259),
    .B(net256),
    .C(_06272_),
    .X(_06283_));
 sky130_fd_sc_hd__a21o_1 _16875_ (.A1(_06270_),
    .A2(_06271_),
    .B1(_05996_),
    .X(_06284_));
 sky130_fd_sc_hd__or4_4 _16876_ (.A(net38),
    .B(net39),
    .C(net40),
    .D(_05477_),
    .X(_06285_));
 sky130_fd_sc_hd__o311a_4 _16877_ (.A1(net39),
    .A2(net40),
    .A3(_05749_),
    .B1(net41),
    .C1(net409),
    .X(_06286_));
 sky130_fd_sc_hd__o211ai_4 _16878_ (.A1(net40),
    .A2(_05989_),
    .B1(net41),
    .C1(net409),
    .Y(_06287_));
 sky130_fd_sc_hd__a21oi_4 _16879_ (.A1(_06285_),
    .A2(net409),
    .B1(net41),
    .Y(_06288_));
 sky130_fd_sc_hd__a21o_4 _16880_ (.A1(_06285_),
    .A2(net409),
    .B1(net41),
    .X(_06290_));
 sky130_fd_sc_hd__a21boi_4 _16881_ (.A1(_06285_),
    .A2(net409),
    .B1_N(net41),
    .Y(_06291_));
 sky130_fd_sc_hd__and3b_4 _16882_ (.A_N(net41),
    .B(_06285_),
    .C(net409),
    .X(_06292_));
 sky130_fd_sc_hd__nor2_8 _16883_ (.A(_06286_),
    .B(_06288_),
    .Y(_06293_));
 sky130_fd_sc_hd__nand2_8 _16884_ (.A(_06287_),
    .B(_06290_),
    .Y(_06294_));
 sky130_fd_sc_hd__a21oi_2 _16885_ (.A1(_06282_),
    .A2(_06283_),
    .B1(_03289_),
    .Y(_06295_));
 sky130_fd_sc_hd__o311ai_2 _16886_ (.A1(_05995_),
    .A2(_06276_),
    .A3(_06279_),
    .B1(_06284_),
    .C1(net1),
    .Y(_06296_));
 sky130_fd_sc_hd__o311a_1 _16887_ (.A1(net259),
    .A2(net256),
    .A3(_06272_),
    .B1(_06282_),
    .C1(_03289_),
    .X(_06297_));
 sky130_fd_sc_hd__o22a_1 _16888_ (.A1(_06291_),
    .A2(_06292_),
    .B1(_06295_),
    .B2(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__a31oi_4 _16889_ (.A1(_06282_),
    .A2(_06283_),
    .A3(_06294_),
    .B1(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__and3_1 _16890_ (.A(_05119_),
    .B(_06003_),
    .C(_06299_),
    .X(_06301_));
 sky130_fd_sc_hd__a21oi_1 _16891_ (.A1(_05119_),
    .A2(_06003_),
    .B1(_06299_),
    .Y(_06302_));
 sky130_fd_sc_hd__nor2_1 _16892_ (.A(_06301_),
    .B(_06302_),
    .Y(net73));
 sky130_fd_sc_hd__o21ai_1 _16893_ (.A1(_06003_),
    .A2(_06299_),
    .B1(_05119_),
    .Y(_06303_));
 sky130_fd_sc_hd__or4_4 _16894_ (.A(net7),
    .B(net8),
    .C(net9),
    .D(_05498_),
    .X(_06304_));
 sky130_fd_sc_hd__and3b_4 _16895_ (.A_N(net10),
    .B(_06304_),
    .C(net410),
    .X(_06305_));
 sky130_fd_sc_hd__inv_4 _16896_ (.A(net284),
    .Y(_06306_));
 sky130_fd_sc_hd__a21boi_4 _16897_ (.A1(_06304_),
    .A2(net410),
    .B1_N(net10),
    .Y(_06307_));
 sky130_fd_sc_hd__a21bo_4 _16898_ (.A1(_06304_),
    .A2(net410),
    .B1_N(net10),
    .X(_06308_));
 sky130_fd_sc_hd__o311a_4 _16899_ (.A1(net8),
    .A2(net9),
    .A3(_05759_),
    .B1(net10),
    .C1(net410),
    .X(_06309_));
 sky130_fd_sc_hd__o211ai_4 _16900_ (.A1(net9),
    .A2(_06008_),
    .B1(net10),
    .C1(net410),
    .Y(_06311_));
 sky130_fd_sc_hd__a21oi_4 _16901_ (.A1(_06304_),
    .A2(net410),
    .B1(net10),
    .Y(_06312_));
 sky130_fd_sc_hd__a21o_4 _16902_ (.A1(_06304_),
    .A2(net410),
    .B1(net10),
    .X(_06313_));
 sky130_fd_sc_hd__nand2_8 _16903_ (.A(_06311_),
    .B(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__nor2_8 _16904_ (.A(_06309_),
    .B(_06312_),
    .Y(_06315_));
 sky130_fd_sc_hd__o32a_1 _16905_ (.A1(_03178_),
    .A2(_06309_),
    .A3(_06312_),
    .B1(net408),
    .B2(_05152_),
    .X(_06316_));
 sky130_fd_sc_hd__a31o_1 _16906_ (.A1(_06313_),
    .A2(net33),
    .A3(_06311_),
    .B1(net405),
    .X(_06317_));
 sky130_fd_sc_hd__o32a_1 _16907_ (.A1(_03178_),
    .A2(_06309_),
    .A3(_06312_),
    .B1(net286),
    .B2(_06012_),
    .X(_06318_));
 sky130_fd_sc_hd__a31o_2 _16908_ (.A1(_06313_),
    .A2(net33),
    .A3(_06311_),
    .B1(net253),
    .X(_06319_));
 sky130_fd_sc_hd__a21oi_2 _16909_ (.A1(_06023_),
    .A2(_06029_),
    .B1(_06024_),
    .Y(_06320_));
 sky130_fd_sc_hd__o21ai_1 _16910_ (.A1(_06030_),
    .A2(_06022_),
    .B1(_06025_),
    .Y(_06322_));
 sky130_fd_sc_hd__and3_1 _16911_ (.A(_06016_),
    .B(_06311_),
    .C(_06313_),
    .X(_06323_));
 sky130_fd_sc_hd__or4_4 _16912_ (.A(_03178_),
    .B(net286),
    .C(_06012_),
    .D(_06314_),
    .X(_06324_));
 sky130_fd_sc_hd__o221ai_4 _16913_ (.A1(_05769_),
    .A2(net254),
    .B1(_06017_),
    .B2(_06314_),
    .C1(_06031_),
    .Y(_06325_));
 sky130_fd_sc_hd__o2111ai_4 _16914_ (.A1(_06017_),
    .A2(_06314_),
    .B1(_06319_),
    .C1(_06025_),
    .D1(_06031_),
    .Y(_06326_));
 sky130_fd_sc_hd__a31o_2 _16915_ (.A1(_06016_),
    .A2(_06311_),
    .A3(_06313_),
    .B1(_06318_),
    .X(_06327_));
 sky130_fd_sc_hd__o2bb2ai_1 _16916_ (.A1_N(_06025_),
    .A2_N(_06031_),
    .B1(_06318_),
    .B2(_06323_),
    .Y(_06328_));
 sky130_fd_sc_hd__a21oi_1 _16917_ (.A1(_06322_),
    .A2(_06327_),
    .B1(_05185_),
    .Y(_06329_));
 sky130_fd_sc_hd__and3_1 _16918_ (.A(_06328_),
    .B(net405),
    .C(_06326_),
    .X(_06330_));
 sky130_fd_sc_hd__nand3_1 _16919_ (.A(_06328_),
    .B(_05174_),
    .C(_06326_),
    .Y(_06331_));
 sky130_fd_sc_hd__a21oi_1 _16920_ (.A1(_06329_),
    .A2(_06326_),
    .B1(_06316_),
    .Y(_06333_));
 sky130_fd_sc_hd__and3_2 _16921_ (.A(_06331_),
    .B(_05392_),
    .C(_06317_),
    .X(_06334_));
 sky130_fd_sc_hd__or4_4 _16922_ (.A(net402),
    .B(net400),
    .C(_06316_),
    .D(_06330_),
    .X(_06335_));
 sky130_fd_sc_hd__or3_1 _16923_ (.A(_05765_),
    .B(net289),
    .C(_06316_),
    .X(_06336_));
 sky130_fd_sc_hd__a21oi_2 _16924_ (.A1(_06329_),
    .A2(_06326_),
    .B1(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__a211o_1 _16925_ (.A1(_06329_),
    .A2(_06326_),
    .B1(_06316_),
    .C1(net262),
    .X(_06338_));
 sky130_fd_sc_hd__a2bb2oi_2 _16926_ (.A1_N(_05765_),
    .A2_N(net289),
    .B1(_06317_),
    .B2(_06331_),
    .Y(_06339_));
 sky130_fd_sc_hd__a2bb2o_1 _16927_ (.A1_N(_05765_),
    .A2_N(net289),
    .B1(_06317_),
    .B2(_06331_),
    .X(_06340_));
 sky130_fd_sc_hd__nor2_2 _16928_ (.A(_06337_),
    .B(_06339_),
    .Y(_06341_));
 sky130_fd_sc_hd__nand3_1 _16929_ (.A(_05531_),
    .B(_05270_),
    .C(_05528_),
    .Y(_06342_));
 sky130_fd_sc_hd__nor3_2 _16930_ (.A(_05788_),
    .B(_06342_),
    .C(_05791_),
    .Y(_06344_));
 sky130_fd_sc_hd__nand4_2 _16931_ (.A(_05792_),
    .B(_05270_),
    .C(_05789_),
    .D(_05532_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand4_4 _16932_ (.A(_06046_),
    .B(_06345_),
    .C(_06040_),
    .D(_06043_),
    .Y(_06346_));
 sky130_fd_sc_hd__a31oi_4 _16933_ (.A1(_06344_),
    .A2(_06040_),
    .A3(_05281_),
    .B1(_06042_),
    .Y(_06347_));
 sky130_fd_sc_hd__nor2_1 _16934_ (.A(_05281_),
    .B(_06345_),
    .Y(_06348_));
 sky130_fd_sc_hd__and3_1 _16935_ (.A(_06348_),
    .B(_06043_),
    .C(_06040_),
    .X(_06349_));
 sky130_fd_sc_hd__nand3_2 _16936_ (.A(_06348_),
    .B(_06043_),
    .C(_06040_),
    .Y(_06350_));
 sky130_fd_sc_hd__a2bb2oi_1 _16937_ (.A1_N(_06034_),
    .A2_N(_06041_),
    .B1(_06040_),
    .B2(_06344_),
    .Y(_06351_));
 sky130_fd_sc_hd__o21a_1 _16938_ (.A1(_06044_),
    .A2(_06047_),
    .B1(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__o21ai_2 _16939_ (.A1(_06044_),
    .A2(_06047_),
    .B1(_06351_),
    .Y(_06353_));
 sky130_fd_sc_hd__nand3_4 _16940_ (.A(_06353_),
    .B(_06341_),
    .C(_06350_),
    .Y(_06355_));
 sky130_fd_sc_hd__o211ai_4 _16941_ (.A1(_06337_),
    .A2(_06339_),
    .B1(_06347_),
    .C1(_06346_),
    .Y(_06356_));
 sky130_fd_sc_hd__o211ai_1 _16942_ (.A1(_06337_),
    .A2(_06339_),
    .B1(_06350_),
    .C1(_06353_),
    .Y(_06357_));
 sky130_fd_sc_hd__o2111ai_2 _16943_ (.A1(_06330_),
    .A2(_06336_),
    .B1(_06340_),
    .C1(_06347_),
    .D1(_06346_),
    .Y(_06358_));
 sky130_fd_sc_hd__a21oi_2 _16944_ (.A1(_06357_),
    .A2(_06358_),
    .B1(_05392_),
    .Y(_06359_));
 sky130_fd_sc_hd__nand3_2 _16945_ (.A(net388),
    .B(_06355_),
    .C(_06356_),
    .Y(_06360_));
 sky130_fd_sc_hd__o22a_4 _16946_ (.A1(_05654_),
    .A2(_05665_),
    .B1(_06334_),
    .B2(_06359_),
    .X(_06361_));
 sky130_fd_sc_hd__a211o_1 _16947_ (.A1(_06335_),
    .A2(_06360_),
    .B1(net384),
    .C1(net383),
    .X(_06362_));
 sky130_fd_sc_hd__a221oi_2 _16948_ (.A1(_05804_),
    .A2(_05806_),
    .B1(_06054_),
    .B2(net293),
    .C1(_05801_),
    .Y(_06363_));
 sky130_fd_sc_hd__a22oi_2 _16949_ (.A1(_06039_),
    .A2(_06057_),
    .B1(_06063_),
    .B2(_06056_),
    .Y(_06364_));
 sky130_fd_sc_hd__o22ai_2 _16950_ (.A1(_06038_),
    .A2(_06058_),
    .B1(_06055_),
    .B2(_06064_),
    .Y(_06366_));
 sky130_fd_sc_hd__a31oi_1 _16951_ (.A1(net388),
    .A2(_06355_),
    .A3(_06356_),
    .B1(net291),
    .Y(_06367_));
 sky130_fd_sc_hd__a311oi_4 _16952_ (.A1(net388),
    .A2(_06355_),
    .A3(_06356_),
    .B1(net291),
    .C1(_06334_),
    .Y(_06368_));
 sky130_fd_sc_hd__nand3_4 _16953_ (.A(_06360_),
    .B(net267),
    .C(_06335_),
    .Y(_06369_));
 sky130_fd_sc_hd__a2bb2oi_2 _16954_ (.A1_N(_05500_),
    .A2_N(_05503_),
    .B1(_06335_),
    .B2(_06360_),
    .Y(_06370_));
 sky130_fd_sc_hd__o22ai_4 _16955_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_06334_),
    .B2(_06359_),
    .Y(_06371_));
 sky130_fd_sc_hd__a21oi_2 _16956_ (.A1(_06335_),
    .A2(_06367_),
    .B1(_06370_),
    .Y(_06372_));
 sky130_fd_sc_hd__nand3_4 _16957_ (.A(_06364_),
    .B(_06369_),
    .C(_06371_),
    .Y(_06373_));
 sky130_fd_sc_hd__o22ai_4 _16958_ (.A1(_06060_),
    .A2(_06363_),
    .B1(_06368_),
    .B2(_06370_),
    .Y(_06374_));
 sky130_fd_sc_hd__o211a_1 _16959_ (.A1(net384),
    .A2(net383),
    .B1(_06373_),
    .C1(_06374_),
    .X(_06375_));
 sky130_fd_sc_hd__o211ai_2 _16960_ (.A1(net384),
    .A2(net383),
    .B1(_06373_),
    .C1(_06374_),
    .Y(_06377_));
 sky130_fd_sc_hd__a31oi_4 _16961_ (.A1(_06373_),
    .A2(_06374_),
    .A3(net359),
    .B1(_06361_),
    .Y(_06378_));
 sky130_fd_sc_hd__a31o_2 _16962_ (.A1(_06373_),
    .A2(_06374_),
    .A3(net359),
    .B1(_06361_),
    .X(_06379_));
 sky130_fd_sc_hd__o21bai_4 _16963_ (.A1(_06082_),
    .A2(_06085_),
    .B1_N(_06077_),
    .Y(_06380_));
 sky130_fd_sc_hd__a311oi_4 _16964_ (.A1(_06373_),
    .A2(_06374_),
    .A3(net359),
    .B1(net293),
    .C1(_06361_),
    .Y(_06381_));
 sky130_fd_sc_hd__a311o_1 _16965_ (.A1(_06373_),
    .A2(_06374_),
    .A3(net359),
    .B1(net293),
    .C1(_06361_),
    .X(_06382_));
 sky130_fd_sc_hd__a2bb2oi_4 _16966_ (.A1_N(_05242_),
    .A2_N(net317),
    .B1(_06362_),
    .B2(_06377_),
    .Y(_06383_));
 sky130_fd_sc_hd__o22ai_4 _16967_ (.A1(_05242_),
    .A2(net317),
    .B1(_06361_),
    .B2(_06375_),
    .Y(_06384_));
 sky130_fd_sc_hd__nand3_4 _16968_ (.A(_06380_),
    .B(_06382_),
    .C(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__o221ai_4 _16969_ (.A1(net299),
    .A2(_06074_),
    .B1(_06381_),
    .B2(_06383_),
    .C1(_06088_),
    .Y(_06386_));
 sky130_fd_sc_hd__and3_2 _16970_ (.A(_06804_),
    .B(_06826_),
    .C(_06379_),
    .X(_06388_));
 sky130_fd_sc_hd__or3_1 _16971_ (.A(net379),
    .B(net378),
    .C(_06378_),
    .X(_06389_));
 sky130_fd_sc_hd__nand3_1 _16972_ (.A(_06385_),
    .B(_06386_),
    .C(net357),
    .Y(_06390_));
 sky130_fd_sc_hd__a31o_1 _16973_ (.A1(_06385_),
    .A2(_06386_),
    .A3(net357),
    .B1(_06388_),
    .X(_06391_));
 sky130_fd_sc_hd__a31oi_4 _16974_ (.A1(_06385_),
    .A2(_06386_),
    .A3(net357),
    .B1(_06388_),
    .Y(_06392_));
 sky130_fd_sc_hd__o311a_2 _16975_ (.A1(net379),
    .A2(net378),
    .A3(_06378_),
    .B1(_06390_),
    .C1(_07724_),
    .X(_06393_));
 sky130_fd_sc_hd__a2bb2oi_2 _16976_ (.A1_N(net339),
    .A2_N(_04184_),
    .B1(_06389_),
    .B2(_06390_),
    .Y(_06394_));
 sky130_fd_sc_hd__a22o_1 _16977_ (.A1(_04173_),
    .A2(_04195_),
    .B1(_06389_),
    .B2(_06390_),
    .X(_06395_));
 sky130_fd_sc_hd__a311oi_4 _16978_ (.A1(_06385_),
    .A2(_06386_),
    .A3(net357),
    .B1(_06388_),
    .C1(net298),
    .Y(_06396_));
 sky130_fd_sc_hd__a311o_1 _16979_ (.A1(_06385_),
    .A2(_06386_),
    .A3(net357),
    .B1(_06388_),
    .C1(net298),
    .X(_06397_));
 sky130_fd_sc_hd__a31o_1 _16980_ (.A1(_05845_),
    .A2(_06099_),
    .A3(_06100_),
    .B1(_06095_),
    .X(_06399_));
 sky130_fd_sc_hd__a31oi_4 _16981_ (.A1(_05845_),
    .A2(_06099_),
    .A3(_06100_),
    .B1(_06095_),
    .Y(_06400_));
 sky130_fd_sc_hd__nand3_2 _16982_ (.A(_06395_),
    .B(_06397_),
    .C(_06400_),
    .Y(_06401_));
 sky130_fd_sc_hd__o21ai_4 _16983_ (.A1(_06394_),
    .A2(_06396_),
    .B1(_06399_),
    .Y(_06402_));
 sky130_fd_sc_hd__o211ai_2 _16984_ (.A1(net373),
    .A2(net371),
    .B1(_06401_),
    .C1(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__or3_1 _16985_ (.A(net373),
    .B(net371),
    .C(_06392_),
    .X(_06404_));
 sky130_fd_sc_hd__o221ai_2 _16986_ (.A1(_06102_),
    .A2(_06098_),
    .B1(_06396_),
    .B2(_06394_),
    .C1(_06096_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand3_1 _16987_ (.A(_06395_),
    .B(_06399_),
    .C(_06397_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand3_2 _16988_ (.A(_06405_),
    .B(_06406_),
    .C(net356),
    .Y(_06407_));
 sky130_fd_sc_hd__o21ai_4 _16989_ (.A1(net355),
    .A2(_06392_),
    .B1(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__a31o_2 _16990_ (.A1(_06402_),
    .A2(net356),
    .A3(_06401_),
    .B1(_06393_),
    .X(_06410_));
 sky130_fd_sc_hd__a311oi_4 _16991_ (.A1(_06401_),
    .A2(_06402_),
    .A3(net356),
    .B1(_02137_),
    .C1(_06393_),
    .Y(_06411_));
 sky130_fd_sc_hd__o211ai_4 _16992_ (.A1(net356),
    .A2(_06391_),
    .B1(_06403_),
    .C1(_02148_),
    .Y(_06412_));
 sky130_fd_sc_hd__a31oi_1 _16993_ (.A1(_06405_),
    .A2(_06406_),
    .A3(net356),
    .B1(_02148_),
    .Y(_06413_));
 sky130_fd_sc_hd__nand3_2 _16994_ (.A(_06407_),
    .B(_02137_),
    .C(_06404_),
    .Y(_06414_));
 sky130_fd_sc_hd__a21oi_2 _16995_ (.A1(_06404_),
    .A2(_06413_),
    .B1(_06411_),
    .Y(_06415_));
 sky130_fd_sc_hd__nand2_1 _16996_ (.A(_06412_),
    .B(_06414_),
    .Y(_06416_));
 sky130_fd_sc_hd__o2111a_1 _16997_ (.A1(_05347_),
    .A2(_05334_),
    .B1(_05346_),
    .C1(_05601_),
    .D1(_05604_),
    .X(_06417_));
 sky130_fd_sc_hd__o2111ai_2 _16998_ (.A1(_05347_),
    .A2(_05334_),
    .B1(_05346_),
    .C1(_05601_),
    .D1(_05604_),
    .Y(_06418_));
 sky130_fd_sc_hd__o21a_1 _16999_ (.A1(_12888_),
    .A2(_05854_),
    .B1(_06417_),
    .X(_06419_));
 sky130_fd_sc_hd__a211oi_2 _17000_ (.A1(_05842_),
    .A2(_05860_),
    .B1(_06418_),
    .C1(_05864_),
    .Y(_06421_));
 sky130_fd_sc_hd__nand3_1 _17001_ (.A(_06419_),
    .B(_06117_),
    .C(_05863_),
    .Y(_06422_));
 sky130_fd_sc_hd__a31oi_1 _17002_ (.A1(_06419_),
    .A2(_06117_),
    .A3(_05863_),
    .B1(_06118_),
    .Y(_06423_));
 sky130_fd_sc_hd__o211ai_4 _17003_ (.A1(_06123_),
    .A2(_06116_),
    .B1(_06119_),
    .C1(_06422_),
    .Y(_06424_));
 sky130_fd_sc_hd__nand4_1 _17004_ (.A(_05863_),
    .B(_06419_),
    .C(_06117_),
    .D(_05350_),
    .Y(_06425_));
 sky130_fd_sc_hd__nand4_4 _17005_ (.A(_06117_),
    .B(_06421_),
    .C(_06119_),
    .D(_05350_),
    .Y(_06426_));
 sky130_fd_sc_hd__a2bb2oi_2 _17006_ (.A1_N(_06118_),
    .A2_N(_06425_),
    .B1(_06127_),
    .B2(_06423_),
    .Y(_06427_));
 sky130_fd_sc_hd__a21oi_2 _17007_ (.A1(_06424_),
    .A2(_06426_),
    .B1(_06416_),
    .Y(_06428_));
 sky130_fd_sc_hd__a21o_1 _17008_ (.A1(_06424_),
    .A2(_06426_),
    .B1(_06416_),
    .X(_06429_));
 sky130_fd_sc_hd__a31oi_2 _17009_ (.A1(_06416_),
    .A2(_06424_),
    .A3(_06426_),
    .B1(_08732_),
    .Y(_06430_));
 sky130_fd_sc_hd__a31o_1 _17010_ (.A1(_06416_),
    .A2(_06424_),
    .A3(_06426_),
    .B1(_08732_),
    .X(_06432_));
 sky130_fd_sc_hd__nand4_4 _17011_ (.A(_06412_),
    .B(_06414_),
    .C(_06424_),
    .D(_06426_),
    .Y(_06433_));
 sky130_fd_sc_hd__a22o_1 _17012_ (.A1(_06412_),
    .A2(_06414_),
    .B1(_06424_),
    .B2(_06426_),
    .X(_06434_));
 sky130_fd_sc_hd__a311o_2 _17013_ (.A1(_06402_),
    .A2(net356),
    .A3(_06401_),
    .B1(net338),
    .C1(_06393_),
    .X(_06435_));
 sky130_fd_sc_hd__o221ai_4 _17014_ (.A1(net353),
    .A2(net352),
    .B1(_06415_),
    .B2(_06427_),
    .C1(_06433_),
    .Y(_06436_));
 sky130_fd_sc_hd__a22oi_4 _17015_ (.A1(_08732_),
    .A2(_06410_),
    .B1(_06430_),
    .B2(_06429_),
    .Y(_06437_));
 sky130_fd_sc_hd__inv_2 _17016_ (.A(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__o221a_2 _17017_ (.A1(net338),
    .A2(_06408_),
    .B1(_06428_),
    .B2(_06432_),
    .C1(_09840_),
    .X(_06439_));
 sky130_fd_sc_hd__a221o_1 _17018_ (.A1(_08732_),
    .A2(_06410_),
    .B1(_06430_),
    .B2(_06429_),
    .C1(net337),
    .X(_06440_));
 sky130_fd_sc_hd__a31oi_2 _17019_ (.A1(_06434_),
    .A2(net338),
    .A3(_06433_),
    .B1(net319),
    .Y(_06441_));
 sky130_fd_sc_hd__and3_2 _17020_ (.A(_06436_),
    .B(net320),
    .C(_06435_),
    .X(_06443_));
 sky130_fd_sc_hd__nand3_2 _17021_ (.A(_06436_),
    .B(net320),
    .C(_06435_),
    .Y(_06444_));
 sky130_fd_sc_hd__o221ai_4 _17022_ (.A1(_08721_),
    .A2(_06408_),
    .B1(_06428_),
    .B2(_06432_),
    .C1(net319),
    .Y(_06445_));
 sky130_fd_sc_hd__o31a_1 _17023_ (.A1(_12867_),
    .A2(_12877_),
    .A3(_06130_),
    .B1(_06135_),
    .X(_06446_));
 sky130_fd_sc_hd__o21ai_1 _17024_ (.A1(_12888_),
    .A2(_06130_),
    .B1(_06135_),
    .Y(_06447_));
 sky130_fd_sc_hd__o21ai_2 _17025_ (.A1(_06137_),
    .A2(_06135_),
    .B1(_06140_),
    .Y(_06448_));
 sky130_fd_sc_hd__o21a_1 _17026_ (.A1(_06137_),
    .A2(_06135_),
    .B1(_06140_),
    .X(_06449_));
 sky130_fd_sc_hd__a21oi_1 _17027_ (.A1(_06444_),
    .A2(_06445_),
    .B1(_06448_),
    .Y(_06450_));
 sky130_fd_sc_hd__o2bb2ai_4 _17028_ (.A1_N(_06444_),
    .A2_N(_06445_),
    .B1(_06446_),
    .B2(_06137_),
    .Y(_06451_));
 sky130_fd_sc_hd__nand3_2 _17029_ (.A(_06444_),
    .B(_06445_),
    .C(_06448_),
    .Y(_06452_));
 sky130_fd_sc_hd__a31o_1 _17030_ (.A1(_06444_),
    .A2(_06445_),
    .A3(_06448_),
    .B1(_09840_),
    .X(_06454_));
 sky130_fd_sc_hd__nand3_1 _17031_ (.A(_06451_),
    .B(_06452_),
    .C(net337),
    .Y(_06455_));
 sky130_fd_sc_hd__a31oi_4 _17032_ (.A1(_06451_),
    .A2(_06452_),
    .A3(net337),
    .B1(_06439_),
    .Y(_06456_));
 sky130_fd_sc_hd__o22ai_4 _17033_ (.A1(net337),
    .A2(_06438_),
    .B1(_06450_),
    .B2(_06454_),
    .Y(_06457_));
 sky130_fd_sc_hd__o22a_1 _17034_ (.A1(net331),
    .A2(_06149_),
    .B1(_06154_),
    .B2(_05892_),
    .X(_06458_));
 sky130_fd_sc_hd__a32oi_4 _17035_ (.A1(net331),
    .A2(_06144_),
    .A3(_06148_),
    .B1(_06155_),
    .B2(_06151_),
    .Y(_06459_));
 sky130_fd_sc_hd__a21boi_1 _17036_ (.A1(_06153_),
    .A2(_06156_),
    .B1_N(_06151_),
    .Y(_06460_));
 sky130_fd_sc_hd__a311oi_4 _17037_ (.A1(_06451_),
    .A2(_06452_),
    .A3(net337),
    .B1(net325),
    .C1(_06439_),
    .Y(_06461_));
 sky130_fd_sc_hd__nand3_2 _17038_ (.A(_06455_),
    .B(_12888_),
    .C(_06440_),
    .Y(_06462_));
 sky130_fd_sc_hd__a2bb2oi_2 _17039_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_06440_),
    .B2(_06455_),
    .Y(_06463_));
 sky130_fd_sc_hd__o21ai_1 _17040_ (.A1(_12845_),
    .A2(_12856_),
    .B1(_06457_),
    .Y(_06465_));
 sky130_fd_sc_hd__o211ai_1 _17041_ (.A1(_06152_),
    .A2(_06458_),
    .B1(_06462_),
    .C1(_06465_),
    .Y(_06466_));
 sky130_fd_sc_hd__o21ai_1 _17042_ (.A1(_06461_),
    .A2(_06463_),
    .B1(_06459_),
    .Y(_06467_));
 sky130_fd_sc_hd__o211ai_2 _17043_ (.A1(net347),
    .A2(net346),
    .B1(_06466_),
    .C1(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__or3_2 _17044_ (.A(net347),
    .B(net346),
    .C(_06456_),
    .X(_06469_));
 sky130_fd_sc_hd__o21ai_1 _17045_ (.A1(_12888_),
    .A2(_06456_),
    .B1(_06459_),
    .Y(_06470_));
 sky130_fd_sc_hd__o22ai_2 _17046_ (.A1(_06152_),
    .A2(_06458_),
    .B1(_06461_),
    .B2(_06463_),
    .Y(_06471_));
 sky130_fd_sc_hd__o221ai_4 _17047_ (.A1(net347),
    .A2(net346),
    .B1(_06461_),
    .B2(_06470_),
    .C1(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__o21ai_2 _17048_ (.A1(net334),
    .A2(_06456_),
    .B1(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__o311a_2 _17049_ (.A1(net347),
    .A2(net346),
    .A3(_06456_),
    .B1(_06472_),
    .C1(_12703_),
    .X(_06474_));
 sky130_fd_sc_hd__a2bb2oi_4 _17050_ (.A1_N(_11210_),
    .A2_N(_11232_),
    .B1(_06469_),
    .B2(_06472_),
    .Y(_06476_));
 sky130_fd_sc_hd__o211ai_4 _17051_ (.A1(_06457_),
    .A2(net334),
    .B1(net330),
    .C1(_06468_),
    .Y(_06477_));
 sky130_fd_sc_hd__o211a_2 _17052_ (.A1(net334),
    .A2(_06456_),
    .B1(net331),
    .C1(_06472_),
    .X(_06478_));
 sky130_fd_sc_hd__o211ai_4 _17053_ (.A1(net334),
    .A2(_06456_),
    .B1(net331),
    .C1(_06472_),
    .Y(_06479_));
 sky130_fd_sc_hd__o21ai_2 _17054_ (.A1(_06172_),
    .A2(_06174_),
    .B1(_06170_),
    .Y(_06480_));
 sky130_fd_sc_hd__o22ai_2 _17055_ (.A1(_06163_),
    .A2(_06171_),
    .B1(_06168_),
    .B2(_06175_),
    .Y(_06481_));
 sky130_fd_sc_hd__nand3_4 _17056_ (.A(_06477_),
    .B(_06479_),
    .C(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__o22ai_4 _17057_ (.A1(_06168_),
    .A2(_06177_),
    .B1(_06476_),
    .B2(_06478_),
    .Y(_06483_));
 sky130_fd_sc_hd__o211ai_2 _17058_ (.A1(net328),
    .A2(_12681_),
    .B1(_06482_),
    .C1(_06483_),
    .Y(_06484_));
 sky130_fd_sc_hd__o211a_1 _17059_ (.A1(_06457_),
    .A2(net334),
    .B1(_12703_),
    .C1(_06468_),
    .X(_06485_));
 sky130_fd_sc_hd__a211o_1 _17060_ (.A1(_06469_),
    .A2(_06472_),
    .B1(net328),
    .C1(_12681_),
    .X(_06487_));
 sky130_fd_sc_hd__a21oi_1 _17061_ (.A1(_06477_),
    .A2(_06479_),
    .B1(_06480_),
    .Y(_06488_));
 sky130_fd_sc_hd__o21ai_1 _17062_ (.A1(_06476_),
    .A2(_06478_),
    .B1(_06481_),
    .Y(_06489_));
 sky130_fd_sc_hd__nand3_2 _17063_ (.A(_06477_),
    .B(_06479_),
    .C(_06480_),
    .Y(_06490_));
 sky130_fd_sc_hd__a31o_1 _17064_ (.A1(_06477_),
    .A2(_06480_),
    .A3(_06479_),
    .B1(_12703_),
    .X(_06491_));
 sky130_fd_sc_hd__a31oi_4 _17065_ (.A1(_06483_),
    .A2(net313),
    .A3(_06482_),
    .B1(_06474_),
    .Y(_06492_));
 sky130_fd_sc_hd__and3_2 _17066_ (.A(_06492_),
    .B(_00044_),
    .C(_00022_),
    .X(_06493_));
 sky130_fd_sc_hd__a311o_2 _17067_ (.A1(_06483_),
    .A2(net313),
    .A3(_06482_),
    .B1(net310),
    .C1(_06474_),
    .X(_06494_));
 sky130_fd_sc_hd__a311oi_4 _17068_ (.A1(_06483_),
    .A2(net313),
    .A3(_06482_),
    .B1(_06474_),
    .C1(_10015_),
    .Y(_06495_));
 sky130_fd_sc_hd__o211ai_4 _17069_ (.A1(net313),
    .A2(_06473_),
    .B1(_06484_),
    .C1(net348),
    .Y(_06496_));
 sky130_fd_sc_hd__a311oi_4 _17070_ (.A1(_06489_),
    .A2(_06490_),
    .A3(net313),
    .B1(_06485_),
    .C1(net348),
    .Y(_06498_));
 sky130_fd_sc_hd__o211ai_4 _17071_ (.A1(_06488_),
    .A2(_06491_),
    .B1(_10015_),
    .C1(_06487_),
    .Y(_06499_));
 sky130_fd_sc_hd__a21oi_2 _17072_ (.A1(_05921_),
    .A2(_05922_),
    .B1(_06187_),
    .Y(_06500_));
 sky130_fd_sc_hd__o31a_4 _17073_ (.A1(_05918_),
    .A2(_06005_),
    .A3(_06187_),
    .B1(_06190_),
    .X(_06501_));
 sky130_fd_sc_hd__o21ai_1 _17074_ (.A1(_06007_),
    .A2(_06187_),
    .B1(_06190_),
    .Y(_06502_));
 sky130_fd_sc_hd__o2111ai_1 _17075_ (.A1(_06007_),
    .A2(_06187_),
    .B1(_06190_),
    .C1(_06496_),
    .D1(_06499_),
    .Y(_06503_));
 sky130_fd_sc_hd__o2bb2ai_1 _17076_ (.A1_N(_06496_),
    .A2_N(_06499_),
    .B1(_06500_),
    .B2(_06189_),
    .Y(_06504_));
 sky130_fd_sc_hd__o21ai_4 _17077_ (.A1(_06495_),
    .A2(_06498_),
    .B1(_06501_),
    .Y(_06505_));
 sky130_fd_sc_hd__o21ai_2 _17078_ (.A1(_06189_),
    .A2(_06500_),
    .B1(_06499_),
    .Y(_06506_));
 sky130_fd_sc_hd__o221ai_4 _17079_ (.A1(_06189_),
    .A2(_06500_),
    .B1(net348),
    .B2(_06492_),
    .C1(_06496_),
    .Y(_06507_));
 sky130_fd_sc_hd__a2bb2oi_2 _17080_ (.A1_N(net324),
    .A2_N(net322),
    .B1(_06503_),
    .B2(_06504_),
    .Y(_06509_));
 sky130_fd_sc_hd__o221ai_4 _17081_ (.A1(net324),
    .A2(net322),
    .B1(_06495_),
    .B2(_06506_),
    .C1(_06505_),
    .Y(_06510_));
 sky130_fd_sc_hd__a31o_1 _17082_ (.A1(_06505_),
    .A2(_06507_),
    .A3(net310),
    .B1(_06493_),
    .X(_06511_));
 sky130_fd_sc_hd__a211o_2 _17083_ (.A1(_06494_),
    .A2(_06510_),
    .B1(net306),
    .C1(net303),
    .X(_06512_));
 sky130_fd_sc_hd__a31o_1 _17084_ (.A1(_06505_),
    .A2(_06507_),
    .A3(net310),
    .B1(_08918_),
    .X(_06513_));
 sky130_fd_sc_hd__a311oi_4 _17085_ (.A1(_06505_),
    .A2(_06507_),
    .A3(net310),
    .B1(_06493_),
    .C1(_08918_),
    .Y(_06514_));
 sky130_fd_sc_hd__o211ai_2 _17086_ (.A1(_08863_),
    .A2(net366),
    .B1(_06494_),
    .C1(_06510_),
    .Y(_06515_));
 sky130_fd_sc_hd__a2bb2oi_1 _17087_ (.A1_N(_08819_),
    .A2_N(net367),
    .B1(_06494_),
    .B2(_06510_),
    .Y(_06516_));
 sky130_fd_sc_hd__o22ai_4 _17088_ (.A1(_08819_),
    .A2(net367),
    .B1(_06493_),
    .B2(_06509_),
    .Y(_06517_));
 sky130_fd_sc_hd__a21oi_1 _17089_ (.A1(_07899_),
    .A2(_06197_),
    .B1(_06200_),
    .Y(_06518_));
 sky130_fd_sc_hd__o32a_1 _17090_ (.A1(net389),
    .A2(net370),
    .A3(_06197_),
    .B1(_06200_),
    .B2(_06203_),
    .X(_06520_));
 sky130_fd_sc_hd__a21oi_2 _17091_ (.A1(_06200_),
    .A2(_06202_),
    .B1(_06203_),
    .Y(_06521_));
 sky130_fd_sc_hd__o22ai_1 _17092_ (.A1(_06203_),
    .A2(_06209_),
    .B1(_06514_),
    .B2(_06516_),
    .Y(_06522_));
 sky130_fd_sc_hd__o221ai_2 _17093_ (.A1(_06201_),
    .A2(_06518_),
    .B1(_06493_),
    .B2(_06513_),
    .C1(_06517_),
    .Y(_06523_));
 sky130_fd_sc_hd__o21ai_1 _17094_ (.A1(_06514_),
    .A2(_06516_),
    .B1(_06521_),
    .Y(_06524_));
 sky130_fd_sc_hd__o211ai_1 _17095_ (.A1(_06203_),
    .A2(_06209_),
    .B1(_06515_),
    .C1(_06517_),
    .Y(_06525_));
 sky130_fd_sc_hd__nand3_2 _17096_ (.A(_06524_),
    .B(_06525_),
    .C(_01962_),
    .Y(_06526_));
 sky130_fd_sc_hd__nand3_2 _17097_ (.A(_06522_),
    .B(_06523_),
    .C(_01962_),
    .Y(_06527_));
 sky130_fd_sc_hd__o31a_1 _17098_ (.A1(_01962_),
    .A2(_06493_),
    .A3(_06509_),
    .B1(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__o311a_2 _17099_ (.A1(_01962_),
    .A2(_06493_),
    .A3(_06509_),
    .B1(_06527_),
    .C1(_07899_),
    .X(_06529_));
 sky130_fd_sc_hd__o211ai_4 _17100_ (.A1(_06511_),
    .A2(_01962_),
    .B1(_07899_),
    .C1(_06527_),
    .Y(_06531_));
 sky130_fd_sc_hd__o211ai_4 _17101_ (.A1(net369),
    .A2(_07866_),
    .B1(_06512_),
    .C1(_06526_),
    .Y(_06532_));
 sky130_fd_sc_hd__o311a_1 _17102_ (.A1(_06332_),
    .A2(_05927_),
    .A3(_05937_),
    .B1(_05948_),
    .C1(_06220_),
    .X(_06533_));
 sky130_fd_sc_hd__o21a_1 _17103_ (.A1(_07044_),
    .A2(_06214_),
    .B1(_06216_),
    .X(_06534_));
 sky130_fd_sc_hd__a21o_1 _17104_ (.A1(_06216_),
    .A2(_06218_),
    .B1(_06219_),
    .X(_06535_));
 sky130_fd_sc_hd__a21oi_1 _17105_ (.A1(_06216_),
    .A2(_06218_),
    .B1(_06219_),
    .Y(_06536_));
 sky130_fd_sc_hd__o2bb2ai_1 _17106_ (.A1_N(_06531_),
    .A2_N(_06532_),
    .B1(_06534_),
    .B2(_06219_),
    .Y(_06537_));
 sky130_fd_sc_hd__o2111ai_1 _17107_ (.A1(_06215_),
    .A2(_06217_),
    .B1(_06220_),
    .C1(_06531_),
    .D1(_06532_),
    .Y(_06538_));
 sky130_fd_sc_hd__o2bb2ai_1 _17108_ (.A1_N(_06531_),
    .A2_N(_06532_),
    .B1(_06533_),
    .B2(_06217_),
    .Y(_06539_));
 sky130_fd_sc_hd__a31oi_2 _17109_ (.A1(_07888_),
    .A2(_06512_),
    .A3(_06526_),
    .B1(_06536_),
    .Y(_06540_));
 sky130_fd_sc_hd__nand3_1 _17110_ (.A(_06531_),
    .B(_06532_),
    .C(_06535_),
    .Y(_06542_));
 sky130_fd_sc_hd__nand3_2 _17111_ (.A(_06539_),
    .B(_06542_),
    .C(net275),
    .Y(_06543_));
 sky130_fd_sc_hd__a211o_1 _17112_ (.A1(_06512_),
    .A2(_06526_),
    .B1(net301),
    .C1(net300),
    .X(_06544_));
 sky130_fd_sc_hd__nand3_1 _17113_ (.A(_06537_),
    .B(_06538_),
    .C(net275),
    .Y(_06545_));
 sky130_fd_sc_hd__nand2_1 _17114_ (.A(_06543_),
    .B(_06544_),
    .Y(_06546_));
 sky130_fd_sc_hd__o21ai_1 _17115_ (.A1(_06332_),
    .A2(_06228_),
    .B1(_06237_),
    .Y(_06547_));
 sky130_fd_sc_hd__nand3_4 _17116_ (.A(_06543_),
    .B(_06544_),
    .C(_07033_),
    .Y(_06548_));
 sky130_fd_sc_hd__o211a_1 _17117_ (.A1(_06528_),
    .A2(net275),
    .B1(_07044_),
    .C1(_06545_),
    .X(_06549_));
 sky130_fd_sc_hd__o211ai_2 _17118_ (.A1(_06528_),
    .A2(net275),
    .B1(_07044_),
    .C1(_06545_),
    .Y(_06550_));
 sky130_fd_sc_hd__o211a_1 _17119_ (.A1(_06229_),
    .A2(_06236_),
    .B1(_06548_),
    .C1(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__o211ai_1 _17120_ (.A1(_06229_),
    .A2(_06236_),
    .B1(_06548_),
    .C1(_06550_),
    .Y(_06553_));
 sky130_fd_sc_hd__a21oi_1 _17121_ (.A1(_06548_),
    .A2(_06550_),
    .B1(_06547_),
    .Y(_06554_));
 sky130_fd_sc_hd__a21o_1 _17122_ (.A1(_06548_),
    .A2(_06550_),
    .B1(_06547_),
    .X(_06555_));
 sky130_fd_sc_hd__o22ai_1 _17123_ (.A1(net297),
    .A2(_05232_),
    .B1(_06551_),
    .B2(_06554_),
    .Y(_06556_));
 sky130_fd_sc_hd__a211o_1 _17124_ (.A1(_06543_),
    .A2(_06544_),
    .B1(net297),
    .C1(_05232_),
    .X(_06557_));
 sky130_fd_sc_hd__o211ai_2 _17125_ (.A1(net297),
    .A2(_05232_),
    .B1(_06553_),
    .C1(_06555_),
    .Y(_06558_));
 sky130_fd_sc_hd__a211o_1 _17126_ (.A1(_06557_),
    .A2(_06558_),
    .B1(_05481_),
    .C1(net269),
    .X(_06559_));
 sky130_fd_sc_hd__a2bb2oi_1 _17127_ (.A1_N(_06245_),
    .A2_N(_06267_),
    .B1(_06557_),
    .B2(_06558_),
    .Y(_06560_));
 sky130_fd_sc_hd__o2111ai_2 _17128_ (.A1(_06546_),
    .A2(net274),
    .B1(_06321_),
    .C1(_06300_),
    .D1(_06556_),
    .Y(_06561_));
 sky130_fd_sc_hd__o211ai_2 _17129_ (.A1(_06289_),
    .A2(net391),
    .B1(_06557_),
    .C1(_06558_),
    .Y(_06562_));
 sky130_fd_sc_hd__o2bb2a_1 _17130_ (.A1_N(_06241_),
    .A2_N(_06255_),
    .B1(_06246_),
    .B2(_06254_),
    .X(_06564_));
 sky130_fd_sc_hd__a21o_1 _17131_ (.A1(_06561_),
    .A2(_06562_),
    .B1(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__nand3_1 _17132_ (.A(_06561_),
    .B(_06562_),
    .C(_06564_),
    .Y(_06566_));
 sky130_fd_sc_hd__nand3_1 _17133_ (.A(_06565_),
    .B(_06566_),
    .C(_05485_),
    .Y(_06567_));
 sky130_fd_sc_hd__a21oi_1 _17134_ (.A1(_06565_),
    .A2(_06566_),
    .B1(_05486_),
    .Y(_06568_));
 sky130_fd_sc_hd__o311a_1 _17135_ (.A1(_05234_),
    .A2(_06551_),
    .A3(_06554_),
    .B1(_06557_),
    .C1(_05486_),
    .X(_06569_));
 sky130_fd_sc_hd__nand2_1 _17136_ (.A(_06559_),
    .B(_06567_),
    .Y(_06570_));
 sky130_fd_sc_hd__o21ai_2 _17137_ (.A1(_06253_),
    .A2(_06262_),
    .B1(_06265_),
    .Y(_06571_));
 sky130_fd_sc_hd__nand4_1 _17138_ (.A(_05982_),
    .B(_05986_),
    .C(_06250_),
    .D(_06252_),
    .Y(_06572_));
 sky130_fd_sc_hd__o211a_1 _17139_ (.A1(net387),
    .A2(_06263_),
    .B1(_06264_),
    .C1(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__a2bb2oi_4 _17140_ (.A1_N(_05763_),
    .A2_N(_05785_),
    .B1(_06264_),
    .B2(_06571_),
    .Y(_06575_));
 sky130_fd_sc_hd__o2111ai_2 _17141_ (.A1(net387),
    .A2(_06263_),
    .B1(_06264_),
    .C1(_05851_),
    .D1(_06572_),
    .Y(_06576_));
 sky130_fd_sc_hd__o21ai_1 _17142_ (.A1(net266),
    .A2(_05751_),
    .B1(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__o21bai_2 _17143_ (.A1(_06575_),
    .A2(_06577_),
    .B1_N(_06570_),
    .Y(_06578_));
 sky130_fd_sc_hd__nand4b_2 _17144_ (.A_N(_06575_),
    .B(net241),
    .C(_06570_),
    .D(_06576_),
    .Y(_06579_));
 sky130_fd_sc_hd__o41a_2 _17145_ (.A1(_06568_),
    .A2(_06569_),
    .A3(_06575_),
    .A4(_06577_),
    .B1(_06578_),
    .X(_06580_));
 sky130_fd_sc_hd__a21boi_2 _17146_ (.A1(_06275_),
    .A2(_05998_),
    .B1_N(_06274_),
    .Y(_06581_));
 sky130_fd_sc_hd__nand3_2 _17147_ (.A(_06281_),
    .B(net387),
    .C(_06274_),
    .Y(_06582_));
 sky130_fd_sc_hd__o211ai_4 _17148_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_06275_),
    .C1(_06277_),
    .Y(_06583_));
 sky130_fd_sc_hd__o2111a_1 _17149_ (.A1(net259),
    .A2(net256),
    .B1(_06582_),
    .C1(_06583_),
    .D1(_06580_),
    .X(_06584_));
 sky130_fd_sc_hd__o2111ai_4 _17150_ (.A1(net259),
    .A2(net256),
    .B1(_06582_),
    .C1(_06583_),
    .D1(_06580_),
    .Y(_06586_));
 sky130_fd_sc_hd__a31oi_2 _17151_ (.A1(_05996_),
    .A2(_06582_),
    .A3(_06583_),
    .B1(_06580_),
    .Y(_06587_));
 sky130_fd_sc_hd__a31o_2 _17152_ (.A1(_05996_),
    .A2(_06582_),
    .A3(_06583_),
    .B1(_06580_),
    .X(_06588_));
 sky130_fd_sc_hd__o211ai_4 _17153_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_06578_),
    .C1(_06579_),
    .Y(_06589_));
 sky130_fd_sc_hd__nand2_1 _17154_ (.A(_06586_),
    .B(_06588_),
    .Y(_06590_));
 sky130_fd_sc_hd__a21oi_2 _17155_ (.A1(_06586_),
    .A2(_06588_),
    .B1(net403),
    .Y(_06591_));
 sky130_fd_sc_hd__o21ai_4 _17156_ (.A1(_06584_),
    .A2(_06587_),
    .B1(_05250_),
    .Y(_06592_));
 sky130_fd_sc_hd__nand3_1 _17157_ (.A(_06588_),
    .B(net403),
    .C(_06586_),
    .Y(_06593_));
 sky130_fd_sc_hd__a31oi_2 _17158_ (.A1(_06588_),
    .A2(net403),
    .A3(_06586_),
    .B1(_06295_),
    .Y(_06594_));
 sky130_fd_sc_hd__a31o_2 _17159_ (.A1(_06588_),
    .A2(net403),
    .A3(_06586_),
    .B1(_06295_),
    .X(_06595_));
 sky130_fd_sc_hd__o41a_1 _17160_ (.A1(net407),
    .A2(_05218_),
    .A3(_06584_),
    .A4(_06587_),
    .B1(_06592_),
    .X(_06597_));
 sky130_fd_sc_hd__a21oi_1 _17161_ (.A1(_06592_),
    .A2(_06593_),
    .B1(_06295_),
    .Y(_06598_));
 sky130_fd_sc_hd__a31o_1 _17162_ (.A1(_06588_),
    .A2(net403),
    .A3(_06586_),
    .B1(_06296_),
    .X(_06599_));
 sky130_fd_sc_hd__o221a_1 _17163_ (.A1(_06591_),
    .A2(_06595_),
    .B1(_06296_),
    .B2(_06597_),
    .C1(net212),
    .X(_06600_));
 sky130_fd_sc_hd__a21oi_1 _17164_ (.A1(_06586_),
    .A2(_06588_),
    .B1(net212),
    .Y(_06601_));
 sky130_fd_sc_hd__o22ai_1 _17165_ (.A1(_06291_),
    .A2(_06292_),
    .B1(_06591_),
    .B2(_06599_),
    .Y(_06602_));
 sky130_fd_sc_hd__o22ai_2 _17166_ (.A1(net212),
    .A2(_06590_),
    .B1(_06598_),
    .B2(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__or4_4 _17167_ (.A(net39),
    .B(net40),
    .C(net41),
    .D(_05749_),
    .X(_06604_));
 sky130_fd_sc_hd__o311a_4 _17168_ (.A1(net40),
    .A2(net41),
    .A3(_05989_),
    .B1(net42),
    .C1(net409),
    .X(_06605_));
 sky130_fd_sc_hd__a21oi_4 _17169_ (.A1(_06604_),
    .A2(net409),
    .B1(net42),
    .Y(_06606_));
 sky130_fd_sc_hd__and3b_4 _17170_ (.A_N(net42),
    .B(_06604_),
    .C(net409),
    .X(_06608_));
 sky130_fd_sc_hd__inv_2 _17171_ (.A(net238),
    .Y(_06609_));
 sky130_fd_sc_hd__a21boi_4 _17172_ (.A1(_06604_),
    .A2(net409),
    .B1_N(net42),
    .Y(_06610_));
 sky130_fd_sc_hd__a21bo_4 _17173_ (.A1(_06604_),
    .A2(net409),
    .B1_N(net42),
    .X(_06611_));
 sky130_fd_sc_hd__nor2_8 _17174_ (.A(_06605_),
    .B(_06606_),
    .Y(_06612_));
 sky130_fd_sc_hd__nor2_8 _17175_ (.A(net238),
    .B(net236),
    .Y(_06613_));
 sky130_fd_sc_hd__o32a_1 _17176_ (.A1(_03289_),
    .A2(_06605_),
    .A3(_06606_),
    .B1(_06600_),
    .B2(_06601_),
    .X(_06614_));
 sky130_fd_sc_hd__nand2_1 _17177_ (.A(net1),
    .B(_06603_),
    .Y(_06615_));
 sky130_fd_sc_hd__a31oi_2 _17178_ (.A1(net1),
    .A2(_06603_),
    .A3(_06612_),
    .B1(_06614_),
    .Y(_06616_));
 sky130_fd_sc_hd__xnor2_1 _17179_ (.A(_06303_),
    .B(_06616_),
    .Y(net74));
 sky130_fd_sc_hd__o32a_1 _17180_ (.A1(_06003_),
    .A2(_06299_),
    .A3(_06616_),
    .B1(_04942_),
    .B2(_04832_),
    .X(_06618_));
 sky130_fd_sc_hd__a21oi_1 _17181_ (.A1(_06562_),
    .A2(_06564_),
    .B1(_06560_),
    .Y(_06619_));
 sky130_fd_sc_hd__a21o_1 _17182_ (.A1(_06562_),
    .A2(_06564_),
    .B1(_06560_),
    .X(_06620_));
 sky130_fd_sc_hd__o21ai_4 _17183_ (.A1(net10),
    .A2(_06304_),
    .B1(net410),
    .Y(_06621_));
 sky130_fd_sc_hd__nor2_8 _17184_ (.A(net11),
    .B(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__or2_4 _17185_ (.A(net11),
    .B(_06621_),
    .X(_06623_));
 sky130_fd_sc_hd__and2_4 _17186_ (.A(_06621_),
    .B(net11),
    .X(_06624_));
 sky130_fd_sc_hd__nand2_4 _17187_ (.A(_06621_),
    .B(net11),
    .Y(_06625_));
 sky130_fd_sc_hd__o311a_4 _17188_ (.A1(net9),
    .A2(net10),
    .A3(_06008_),
    .B1(net11),
    .C1(net410),
    .X(_06626_));
 sky130_fd_sc_hd__and2b_4 _17189_ (.A_N(net11),
    .B(_06621_),
    .X(_06627_));
 sky130_fd_sc_hd__nor2_8 _17190_ (.A(_06622_),
    .B(_06624_),
    .Y(_06629_));
 sky130_fd_sc_hd__nor2_4 _17191_ (.A(_06626_),
    .B(_06627_),
    .Y(_06630_));
 sky130_fd_sc_hd__o21a_2 _17192_ (.A1(_06622_),
    .A2(_06624_),
    .B1(net33),
    .X(_06631_));
 sky130_fd_sc_hd__or4_4 _17193_ (.A(_06626_),
    .B(_03178_),
    .C(_06314_),
    .D(_06627_),
    .X(_06632_));
 sky130_fd_sc_hd__or3_4 _17194_ (.A(_06305_),
    .B(net283),
    .C(_06631_),
    .X(_06633_));
 sky130_fd_sc_hd__nand2_1 _17195_ (.A(_06632_),
    .B(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__nand4_4 _17196_ (.A(_06319_),
    .B(_06325_),
    .C(_06632_),
    .D(_06633_),
    .Y(_06635_));
 sky130_fd_sc_hd__o211ai_4 _17197_ (.A1(_06327_),
    .A2(_06320_),
    .B1(_06324_),
    .C1(_06634_),
    .Y(_06636_));
 sky130_fd_sc_hd__nand3_1 _17198_ (.A(_06635_),
    .B(_06636_),
    .C(net405),
    .Y(_06637_));
 sky130_fd_sc_hd__o221a_1 _17199_ (.A1(_05130_),
    .A2(_05152_),
    .B1(_06622_),
    .B2(_06624_),
    .C1(net33),
    .X(_06638_));
 sky130_fd_sc_hd__or4_1 _17200_ (.A(_03178_),
    .B(net405),
    .C(_06626_),
    .D(_06627_),
    .X(_06640_));
 sky130_fd_sc_hd__o31a_2 _17201_ (.A1(_03178_),
    .A2(net405),
    .A3(net234),
    .B1(_06637_),
    .X(_06641_));
 sky130_fd_sc_hd__or3_1 _17202_ (.A(net402),
    .B(net400),
    .C(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__a311oi_4 _17203_ (.A1(_06635_),
    .A2(_06636_),
    .A3(net405),
    .B1(_06638_),
    .C1(net253),
    .Y(_06643_));
 sky130_fd_sc_hd__a311o_1 _17204_ (.A1(_06635_),
    .A2(_06636_),
    .A3(net405),
    .B1(_06638_),
    .C1(net253),
    .X(_06644_));
 sky130_fd_sc_hd__a21oi_2 _17205_ (.A1(_06637_),
    .A2(_06640_),
    .B1(net254),
    .Y(_06645_));
 sky130_fd_sc_hd__a21o_1 _17206_ (.A1(_06637_),
    .A2(_06640_),
    .B1(net254),
    .X(_06646_));
 sky130_fd_sc_hd__nor2_2 _17207_ (.A(_06643_),
    .B(_06645_),
    .Y(_06647_));
 sky130_fd_sc_hd__nand3_2 _17208_ (.A(_06338_),
    .B(_06346_),
    .C(_06347_),
    .Y(_06648_));
 sky130_fd_sc_hd__o2111ai_4 _17209_ (.A1(net261),
    .A2(_06333_),
    .B1(_06644_),
    .C1(_06646_),
    .D1(_06648_),
    .Y(_06649_));
 sky130_fd_sc_hd__o211ai_2 _17210_ (.A1(_06643_),
    .A2(_06645_),
    .B1(_06338_),
    .C1(_06355_),
    .Y(_06651_));
 sky130_fd_sc_hd__o211ai_4 _17211_ (.A1(net402),
    .A2(_05370_),
    .B1(_06649_),
    .C1(_06651_),
    .Y(_06652_));
 sky130_fd_sc_hd__o21ai_1 _17212_ (.A1(net388),
    .A2(_06641_),
    .B1(_06652_),
    .Y(_06653_));
 sky130_fd_sc_hd__inv_2 _17213_ (.A(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__and3_2 _17214_ (.A(_05687_),
    .B(_05709_),
    .C(_06653_),
    .X(_06655_));
 sky130_fd_sc_hd__a211o_1 _17215_ (.A1(_06642_),
    .A2(_06652_),
    .B1(net384),
    .C1(net383),
    .X(_06656_));
 sky130_fd_sc_hd__a2bb2oi_2 _17216_ (.A1_N(_05760_),
    .A2_N(net290),
    .B1(_06642_),
    .B2(_06652_),
    .Y(_06657_));
 sky130_fd_sc_hd__a22o_1 _17217_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_06642_),
    .B2(_06652_),
    .X(_06658_));
 sky130_fd_sc_hd__o211a_1 _17218_ (.A1(net388),
    .A2(_06641_),
    .B1(net262),
    .C1(_06652_),
    .X(_06659_));
 sky130_fd_sc_hd__o211ai_4 _17219_ (.A1(net388),
    .A2(_06641_),
    .B1(net262),
    .C1(_06652_),
    .Y(_06660_));
 sky130_fd_sc_hd__nor2_2 _17220_ (.A(_06657_),
    .B(_06659_),
    .Y(_06662_));
 sky130_fd_sc_hd__nor4_1 _17221_ (.A(_05550_),
    .B(_05552_),
    .C(_05801_),
    .D(_05803_),
    .Y(_06663_));
 sky130_fd_sc_hd__nand4_2 _17222_ (.A(_05551_),
    .B(_05553_),
    .C(_05802_),
    .D(_05804_),
    .Y(_06664_));
 sky130_fd_sc_hd__nor3_1 _17223_ (.A(_06055_),
    .B(_06060_),
    .C(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__nand3_1 _17224_ (.A(_06369_),
    .B(_06663_),
    .C(_06062_),
    .Y(_06666_));
 sky130_fd_sc_hd__a31oi_2 _17225_ (.A1(_06062_),
    .A2(_06369_),
    .A3(_06663_),
    .B1(_06370_),
    .Y(_06667_));
 sky130_fd_sc_hd__o211ai_4 _17226_ (.A1(_06368_),
    .A2(_06366_),
    .B1(_06666_),
    .C1(_06371_),
    .Y(_06668_));
 sky130_fd_sc_hd__nor4_2 _17227_ (.A(_05548_),
    .B(_06055_),
    .C(_06060_),
    .D(_06664_),
    .Y(_06669_));
 sky130_fd_sc_hd__nand4_4 _17228_ (.A(_06665_),
    .B(_06371_),
    .C(_06369_),
    .D(_05549_),
    .Y(_06670_));
 sky130_fd_sc_hd__a22oi_4 _17229_ (.A1(_06372_),
    .A2(_06669_),
    .B1(_06667_),
    .B2(_06373_),
    .Y(_06671_));
 sky130_fd_sc_hd__a22o_1 _17230_ (.A1(_06372_),
    .A2(_06669_),
    .B1(_06667_),
    .B2(_06373_),
    .X(_06673_));
 sky130_fd_sc_hd__nand4_4 _17231_ (.A(_06658_),
    .B(_06660_),
    .C(_06668_),
    .D(_06670_),
    .Y(_06674_));
 sky130_fd_sc_hd__a22o_1 _17232_ (.A1(_06658_),
    .A2(_06660_),
    .B1(_06668_),
    .B2(_06670_),
    .X(_06675_));
 sky130_fd_sc_hd__o221a_1 _17233_ (.A1(net384),
    .A2(net383),
    .B1(_06662_),
    .B2(_06671_),
    .C1(_06674_),
    .X(_06676_));
 sky130_fd_sc_hd__o221ai_4 _17234_ (.A1(net384),
    .A2(net383),
    .B1(_06662_),
    .B2(_06671_),
    .C1(_06674_),
    .Y(_06677_));
 sky130_fd_sc_hd__o211a_1 _17235_ (.A1(_06655_),
    .A2(_06676_),
    .B1(_06804_),
    .C1(_06826_),
    .X(_06678_));
 sky130_fd_sc_hd__a211o_2 _17236_ (.A1(_06656_),
    .A2(_06677_),
    .B1(net379),
    .C1(net378),
    .X(_06679_));
 sky130_fd_sc_hd__o221a_1 _17237_ (.A1(net295),
    .A2(_06378_),
    .B1(_06084_),
    .B2(_06085_),
    .C1(_06078_),
    .X(_06680_));
 sky130_fd_sc_hd__o221ai_4 _17238_ (.A1(net295),
    .A2(_06378_),
    .B1(_06084_),
    .B2(_06085_),
    .C1(_06078_),
    .Y(_06681_));
 sky130_fd_sc_hd__o32ai_4 _17239_ (.A1(_05242_),
    .A2(net314),
    .A3(_06379_),
    .B1(_06383_),
    .B2(_06380_),
    .Y(_06682_));
 sky130_fd_sc_hd__a311oi_4 _17240_ (.A1(_06675_),
    .A2(net359),
    .A3(_06674_),
    .B1(net291),
    .C1(_06655_),
    .Y(_06684_));
 sky130_fd_sc_hd__o211ai_4 _17241_ (.A1(net359),
    .A2(_06654_),
    .B1(net267),
    .C1(_06677_),
    .Y(_06685_));
 sky130_fd_sc_hd__a2bb2oi_4 _17242_ (.A1_N(_05500_),
    .A2_N(_05503_),
    .B1(_06656_),
    .B2(_06677_),
    .Y(_06686_));
 sky130_fd_sc_hd__o22ai_4 _17243_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_06655_),
    .B2(_06676_),
    .Y(_06687_));
 sky130_fd_sc_hd__o2111ai_4 _17244_ (.A1(net293),
    .A2(_06379_),
    .B1(_06681_),
    .C1(_06685_),
    .D1(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__o22ai_4 _17245_ (.A1(_06381_),
    .A2(_06680_),
    .B1(_06684_),
    .B2(_06686_),
    .Y(_06689_));
 sky130_fd_sc_hd__o211ai_4 _17246_ (.A1(net379),
    .A2(net378),
    .B1(_06688_),
    .C1(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__a31o_2 _17247_ (.A1(_06688_),
    .A2(_06689_),
    .A3(net357),
    .B1(_06678_),
    .X(_06691_));
 sky130_fd_sc_hd__o221a_1 _17248_ (.A1(_06102_),
    .A2(_06098_),
    .B1(net299),
    .B2(_06392_),
    .C1(_06096_),
    .X(_06692_));
 sky130_fd_sc_hd__nor2_1 _17249_ (.A(_06396_),
    .B(_06400_),
    .Y(_06693_));
 sky130_fd_sc_hd__o21ai_2 _17250_ (.A1(_06396_),
    .A2(_06400_),
    .B1(_06395_),
    .Y(_06695_));
 sky130_fd_sc_hd__a311oi_4 _17251_ (.A1(_06688_),
    .A2(_06689_),
    .A3(net357),
    .B1(net293),
    .C1(_06678_),
    .Y(_06696_));
 sky130_fd_sc_hd__o211ai_4 _17252_ (.A1(_05246_),
    .A2(_05247_),
    .B1(_06679_),
    .C1(_06690_),
    .Y(_06697_));
 sky130_fd_sc_hd__a2bb2oi_2 _17253_ (.A1_N(_05242_),
    .A2_N(net314),
    .B1(_06679_),
    .B2(_06690_),
    .Y(_06698_));
 sky130_fd_sc_hd__a22o_1 _17254_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_06679_),
    .B2(_06690_),
    .X(_06699_));
 sky130_fd_sc_hd__o211ai_2 _17255_ (.A1(_06396_),
    .A2(_06692_),
    .B1(_06697_),
    .C1(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__o22ai_2 _17256_ (.A1(_06394_),
    .A2(_06693_),
    .B1(_06696_),
    .B2(_06698_),
    .Y(_06701_));
 sky130_fd_sc_hd__nand3_4 _17257_ (.A(_06700_),
    .B(_06701_),
    .C(net356),
    .Y(_06702_));
 sky130_fd_sc_hd__a211o_1 _17258_ (.A1(_06679_),
    .A2(_06690_),
    .B1(net373),
    .C1(net371),
    .X(_06703_));
 sky130_fd_sc_hd__nand3_1 _17259_ (.A(_06699_),
    .B(_06695_),
    .C(_06697_),
    .Y(_06704_));
 sky130_fd_sc_hd__o22ai_1 _17260_ (.A1(_06396_),
    .A2(_06692_),
    .B1(_06696_),
    .B2(_06698_),
    .Y(_06706_));
 sky130_fd_sc_hd__nand3_1 _17261_ (.A(_06704_),
    .B(_06706_),
    .C(net356),
    .Y(_06707_));
 sky130_fd_sc_hd__o21ai_4 _17262_ (.A1(net355),
    .A2(_06691_),
    .B1(_06702_),
    .Y(_06708_));
 sky130_fd_sc_hd__o211ai_4 _17263_ (.A1(_06691_),
    .A2(net355),
    .B1(net298),
    .C1(_06702_),
    .Y(_06709_));
 sky130_fd_sc_hd__nand3_2 _17264_ (.A(_06707_),
    .B(net299),
    .C(_06703_),
    .Y(_06710_));
 sky130_fd_sc_hd__nand2_1 _17265_ (.A(_06709_),
    .B(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__a21oi_4 _17266_ (.A1(_06424_),
    .A2(_06426_),
    .B1(_06411_),
    .Y(_06712_));
 sky130_fd_sc_hd__o211ai_4 _17267_ (.A1(_06408_),
    .A2(_02148_),
    .B1(_06710_),
    .C1(_06709_),
    .Y(_06713_));
 sky130_fd_sc_hd__o211a_1 _17268_ (.A1(_02137_),
    .A2(_06410_),
    .B1(_06433_),
    .C1(_06711_),
    .X(_06714_));
 sky130_fd_sc_hd__o211ai_2 _17269_ (.A1(_02137_),
    .A2(_06410_),
    .B1(_06433_),
    .C1(_06711_),
    .Y(_06715_));
 sky130_fd_sc_hd__o211a_4 _17270_ (.A1(_06691_),
    .A2(net355),
    .B1(_08732_),
    .C1(_06702_),
    .X(_06717_));
 sky130_fd_sc_hd__inv_2 _17271_ (.A(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__o22ai_2 _17272_ (.A1(net353),
    .A2(net352),
    .B1(_06712_),
    .B2(_06713_),
    .Y(_06719_));
 sky130_fd_sc_hd__o211ai_4 _17273_ (.A1(_06712_),
    .A2(_06713_),
    .B1(net338),
    .C1(_06715_),
    .Y(_06720_));
 sky130_fd_sc_hd__o22ai_4 _17274_ (.A1(net338),
    .A2(_06708_),
    .B1(_06719_),
    .B2(_06714_),
    .Y(_06721_));
 sky130_fd_sc_hd__or3_1 _17275_ (.A(net350),
    .B(net349),
    .C(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__a22oi_4 _17276_ (.A1(_06138_),
    .A2(_06447_),
    .B1(_06437_),
    .B2(net319),
    .Y(_06723_));
 sky130_fd_sc_hd__a22oi_4 _17277_ (.A1(_06435_),
    .A2(_06441_),
    .B1(_06445_),
    .B2(_06449_),
    .Y(_06724_));
 sky130_fd_sc_hd__a2bb2oi_4 _17278_ (.A1_N(_02049_),
    .A2_N(net342),
    .B1(_06718_),
    .B2(_06720_),
    .Y(_06725_));
 sky130_fd_sc_hd__o21ai_2 _17279_ (.A1(_02049_),
    .A2(net342),
    .B1(_06721_),
    .Y(_06726_));
 sky130_fd_sc_hd__o21ai_4 _17280_ (.A1(_02093_),
    .A2(_02115_),
    .B1(_06720_),
    .Y(_06728_));
 sky130_fd_sc_hd__o221a_1 _17281_ (.A1(net338),
    .A2(_06708_),
    .B1(_06719_),
    .B2(_06714_),
    .C1(_02137_),
    .X(_06729_));
 sky130_fd_sc_hd__o21a_1 _17282_ (.A1(_06717_),
    .A2(_06728_),
    .B1(_06726_),
    .X(_06730_));
 sky130_fd_sc_hd__o211ai_4 _17283_ (.A1(_06717_),
    .A2(_06728_),
    .B1(_06724_),
    .C1(_06726_),
    .Y(_06731_));
 sky130_fd_sc_hd__o22ai_4 _17284_ (.A1(_06443_),
    .A2(_06723_),
    .B1(_06725_),
    .B2(_06729_),
    .Y(_06732_));
 sky130_fd_sc_hd__o21ai_1 _17285_ (.A1(_06725_),
    .A2(_06729_),
    .B1(_06724_),
    .Y(_06733_));
 sky130_fd_sc_hd__o221ai_2 _17286_ (.A1(_06443_),
    .A2(_06723_),
    .B1(_06728_),
    .B2(_06717_),
    .C1(_06726_),
    .Y(_06734_));
 sky130_fd_sc_hd__nand3_2 _17287_ (.A(_06733_),
    .B(_06734_),
    .C(net337),
    .Y(_06735_));
 sky130_fd_sc_hd__and3_1 _17288_ (.A(_06721_),
    .B(_09818_),
    .C(_09796_),
    .X(_06736_));
 sky130_fd_sc_hd__a211o_1 _17289_ (.A1(_06718_),
    .A2(_06720_),
    .B1(_09785_),
    .C1(net349),
    .X(_06737_));
 sky130_fd_sc_hd__o211ai_2 _17290_ (.A1(net350),
    .A2(net349),
    .B1(_06731_),
    .C1(_06732_),
    .Y(_06739_));
 sky130_fd_sc_hd__o311a_4 _17291_ (.A1(net350),
    .A2(net349),
    .A3(_06721_),
    .B1(_06735_),
    .C1(_11079_),
    .X(_06740_));
 sky130_fd_sc_hd__inv_2 _17292_ (.A(_06740_),
    .Y(_06741_));
 sky130_fd_sc_hd__a311oi_4 _17293_ (.A1(_06731_),
    .A2(_06732_),
    .A3(net337),
    .B1(_06736_),
    .C1(net319),
    .Y(_06742_));
 sky130_fd_sc_hd__nand3_4 _17294_ (.A(_06739_),
    .B(net320),
    .C(_06737_),
    .Y(_06743_));
 sky130_fd_sc_hd__o311a_2 _17295_ (.A1(net350),
    .A2(net349),
    .A3(_06721_),
    .B1(_06735_),
    .C1(net319),
    .X(_06744_));
 sky130_fd_sc_hd__o211ai_4 _17296_ (.A1(_00174_),
    .A2(_00196_),
    .B1(_06722_),
    .C1(_06735_),
    .Y(_06745_));
 sky130_fd_sc_hd__o21a_1 _17297_ (.A1(_12888_),
    .A2(_06456_),
    .B1(_06460_),
    .X(_06746_));
 sky130_fd_sc_hd__o21ai_1 _17298_ (.A1(_06460_),
    .A2(_06461_),
    .B1(_06465_),
    .Y(_06747_));
 sky130_fd_sc_hd__a21oi_2 _17299_ (.A1(_06459_),
    .A2(_06462_),
    .B1(_06463_),
    .Y(_06748_));
 sky130_fd_sc_hd__o2bb2ai_4 _17300_ (.A1_N(_06743_),
    .A2_N(_06745_),
    .B1(_06746_),
    .B2(_06461_),
    .Y(_06750_));
 sky130_fd_sc_hd__nand3_4 _17301_ (.A(_06747_),
    .B(_06745_),
    .C(_06743_),
    .Y(_06751_));
 sky130_fd_sc_hd__nand3_1 _17302_ (.A(_06750_),
    .B(_06751_),
    .C(net334),
    .Y(_06752_));
 sky130_fd_sc_hd__a31oi_4 _17303_ (.A1(_06750_),
    .A2(_06751_),
    .A3(net334),
    .B1(_06740_),
    .Y(_06753_));
 sky130_fd_sc_hd__a31o_2 _17304_ (.A1(_06750_),
    .A2(_06751_),
    .A3(net334),
    .B1(_06740_),
    .X(_06754_));
 sky130_fd_sc_hd__a21oi_1 _17305_ (.A1(_06473_),
    .A2(net330),
    .B1(_06480_),
    .Y(_06755_));
 sky130_fd_sc_hd__a32oi_4 _17306_ (.A1(_06472_),
    .A2(net331),
    .A3(_06469_),
    .B1(_06170_),
    .B2(_06178_),
    .Y(_06756_));
 sky130_fd_sc_hd__a311oi_4 _17307_ (.A1(_06750_),
    .A2(_06751_),
    .A3(net334),
    .B1(net325),
    .C1(_06740_),
    .Y(_06757_));
 sky130_fd_sc_hd__a311o_1 _17308_ (.A1(_06750_),
    .A2(_06751_),
    .A3(net334),
    .B1(net325),
    .C1(_06740_),
    .X(_06758_));
 sky130_fd_sc_hd__a2bb2oi_4 _17309_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_06741_),
    .B2(_06752_),
    .Y(_06759_));
 sky130_fd_sc_hd__o21ai_1 _17310_ (.A1(_12845_),
    .A2(_12856_),
    .B1(_06754_),
    .Y(_06761_));
 sky130_fd_sc_hd__o211ai_2 _17311_ (.A1(_06478_),
    .A2(_06755_),
    .B1(_06758_),
    .C1(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__o22ai_2 _17312_ (.A1(_06476_),
    .A2(_06756_),
    .B1(_06757_),
    .B2(_06759_),
    .Y(_06763_));
 sky130_fd_sc_hd__o211ai_2 _17313_ (.A1(_06476_),
    .A2(_06756_),
    .B1(_06758_),
    .C1(_06761_),
    .Y(_06764_));
 sky130_fd_sc_hd__o22ai_2 _17314_ (.A1(_06478_),
    .A2(_06755_),
    .B1(_06757_),
    .B2(_06759_),
    .Y(_06765_));
 sky130_fd_sc_hd__nand3_4 _17315_ (.A(_06762_),
    .B(_06763_),
    .C(net313),
    .Y(_06766_));
 sky130_fd_sc_hd__a21oi_1 _17316_ (.A1(_06741_),
    .A2(_06752_),
    .B1(net313),
    .Y(_06767_));
 sky130_fd_sc_hd__inv_2 _17317_ (.A(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__nand3_2 _17318_ (.A(_06764_),
    .B(_06765_),
    .C(net312),
    .Y(_06769_));
 sky130_fd_sc_hd__o21ai_4 _17319_ (.A1(net313),
    .A2(_06754_),
    .B1(_06766_),
    .Y(_06770_));
 sky130_fd_sc_hd__a311o_2 _17320_ (.A1(_06764_),
    .A2(_06765_),
    .A3(net312),
    .B1(_06767_),
    .C1(net310),
    .X(_06772_));
 sky130_fd_sc_hd__o211a_2 _17321_ (.A1(net313),
    .A2(_06753_),
    .B1(net331),
    .C1(_06769_),
    .X(_06773_));
 sky130_fd_sc_hd__o211ai_4 _17322_ (.A1(net313),
    .A2(_06753_),
    .B1(net331),
    .C1(_06769_),
    .Y(_06774_));
 sky130_fd_sc_hd__o211a_1 _17323_ (.A1(_06754_),
    .A2(net313),
    .B1(net330),
    .C1(_06766_),
    .X(_06775_));
 sky130_fd_sc_hd__o211ai_4 _17324_ (.A1(_06754_),
    .A2(net313),
    .B1(net330),
    .C1(_06766_),
    .Y(_06776_));
 sky130_fd_sc_hd__a21oi_1 _17325_ (.A1(_06492_),
    .A2(net348),
    .B1(_06502_),
    .Y(_06777_));
 sky130_fd_sc_hd__a31o_1 _17326_ (.A1(_06492_),
    .A2(_10004_),
    .A3(_09982_),
    .B1(_06502_),
    .X(_06778_));
 sky130_fd_sc_hd__a21oi_1 _17327_ (.A1(_06499_),
    .A2(_06502_),
    .B1(_06495_),
    .Y(_06779_));
 sky130_fd_sc_hd__o2111ai_1 _17328_ (.A1(_06498_),
    .A2(_06501_),
    .B1(_06774_),
    .C1(_06776_),
    .D1(_06496_),
    .Y(_06780_));
 sky130_fd_sc_hd__a22o_1 _17329_ (.A1(_06496_),
    .A2(_06506_),
    .B1(_06774_),
    .B2(_06776_),
    .X(_06781_));
 sky130_fd_sc_hd__o211ai_2 _17330_ (.A1(net324),
    .A2(net322),
    .B1(_06780_),
    .C1(_06781_),
    .Y(_06783_));
 sky130_fd_sc_hd__a211o_1 _17331_ (.A1(_06768_),
    .A2(_06769_),
    .B1(net324),
    .C1(_00033_),
    .X(_06784_));
 sky130_fd_sc_hd__o2bb2ai_1 _17332_ (.A1_N(_06774_),
    .A2_N(_06776_),
    .B1(_06777_),
    .B2(_06498_),
    .Y(_06785_));
 sky130_fd_sc_hd__o2111ai_4 _17333_ (.A1(net348),
    .A2(_06492_),
    .B1(_06774_),
    .C1(_06776_),
    .D1(_06778_),
    .Y(_06786_));
 sky130_fd_sc_hd__nand3_4 _17334_ (.A(_06785_),
    .B(_06786_),
    .C(net310),
    .Y(_06787_));
 sky130_fd_sc_hd__o21ai_2 _17335_ (.A1(net310),
    .A2(_06770_),
    .B1(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__a2bb2oi_2 _17336_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_06784_),
    .B2(_06787_),
    .Y(_06789_));
 sky130_fd_sc_hd__nand4_4 _17337_ (.A(_09982_),
    .B(_10004_),
    .C(_06772_),
    .D(_06783_),
    .Y(_06790_));
 sky130_fd_sc_hd__o221a_2 _17338_ (.A1(_09971_),
    .A2(net363),
    .B1(net310),
    .B2(_06770_),
    .C1(_06787_),
    .X(_06791_));
 sky130_fd_sc_hd__o221ai_4 _17339_ (.A1(_09971_),
    .A2(net363),
    .B1(net310),
    .B2(_06770_),
    .C1(_06787_),
    .Y(_06792_));
 sky130_fd_sc_hd__a21oi_2 _17340_ (.A1(_06520_),
    .A2(_06515_),
    .B1(_06516_),
    .Y(_06794_));
 sky130_fd_sc_hd__o21ai_2 _17341_ (.A1(_06521_),
    .A2(_06514_),
    .B1(_06517_),
    .Y(_06795_));
 sky130_fd_sc_hd__o21ai_4 _17342_ (.A1(_06789_),
    .A2(_06791_),
    .B1(_06794_),
    .Y(_06796_));
 sky130_fd_sc_hd__nand3_4 _17343_ (.A(_06790_),
    .B(_06792_),
    .C(_06795_),
    .Y(_06797_));
 sky130_fd_sc_hd__o2111ai_4 _17344_ (.A1(_06521_),
    .A2(_06514_),
    .B1(_06517_),
    .C1(_06790_),
    .D1(_06792_),
    .Y(_06798_));
 sky130_fd_sc_hd__o21ai_1 _17345_ (.A1(_06789_),
    .A2(_06791_),
    .B1(_06795_),
    .Y(_06799_));
 sky130_fd_sc_hd__o211ai_4 _17346_ (.A1(net306),
    .A2(net303),
    .B1(_06798_),
    .C1(_06799_),
    .Y(_06800_));
 sky130_fd_sc_hd__and3_2 _17347_ (.A(_01973_),
    .B(_06772_),
    .C(_06783_),
    .X(_06801_));
 sky130_fd_sc_hd__a211o_1 _17348_ (.A1(_06784_),
    .A2(_06787_),
    .B1(net306),
    .C1(net303),
    .X(_06802_));
 sky130_fd_sc_hd__nand3_2 _17349_ (.A(_06796_),
    .B(_06797_),
    .C(_01962_),
    .Y(_06803_));
 sky130_fd_sc_hd__a31oi_4 _17350_ (.A1(_06796_),
    .A2(_06797_),
    .A3(_01962_),
    .B1(_06801_),
    .Y(_06805_));
 sky130_fd_sc_hd__o221a_2 _17351_ (.A1(_03986_),
    .A2(_03997_),
    .B1(_06788_),
    .B2(net280),
    .C1(_06800_),
    .X(_06806_));
 sky130_fd_sc_hd__or3_1 _17352_ (.A(net301),
    .B(net300),
    .C(_06805_),
    .X(_06807_));
 sky130_fd_sc_hd__a21oi_2 _17353_ (.A1(_06532_),
    .A2(_06535_),
    .B1(_06529_),
    .Y(_06808_));
 sky130_fd_sc_hd__a311oi_4 _17354_ (.A1(_06796_),
    .A2(_06797_),
    .A3(_01962_),
    .B1(_06801_),
    .C1(_08918_),
    .Y(_06809_));
 sky130_fd_sc_hd__o211ai_2 _17355_ (.A1(_08863_),
    .A2(net366),
    .B1(_06802_),
    .C1(_06803_),
    .Y(_06810_));
 sky130_fd_sc_hd__a2bb2oi_1 _17356_ (.A1_N(_08819_),
    .A2_N(net367),
    .B1(_06802_),
    .B2(_06803_),
    .Y(_06811_));
 sky130_fd_sc_hd__o211ai_4 _17357_ (.A1(net280),
    .A2(_06788_),
    .B1(_06800_),
    .C1(_08918_),
    .Y(_06812_));
 sky130_fd_sc_hd__nand3_1 _17358_ (.A(_06808_),
    .B(_06810_),
    .C(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__o22ai_1 _17359_ (.A1(_06529_),
    .A2(_06540_),
    .B1(_06809_),
    .B2(_06811_),
    .Y(_06814_));
 sky130_fd_sc_hd__o211ai_4 _17360_ (.A1(_06529_),
    .A2(_06540_),
    .B1(_06810_),
    .C1(_06812_),
    .Y(_06816_));
 sky130_fd_sc_hd__o21ai_2 _17361_ (.A1(_06809_),
    .A2(_06811_),
    .B1(_06808_),
    .Y(_06817_));
 sky130_fd_sc_hd__a2bb2oi_2 _17362_ (.A1_N(net301),
    .A2_N(net300),
    .B1(_06813_),
    .B2(_06814_),
    .Y(_06818_));
 sky130_fd_sc_hd__nand3_2 _17363_ (.A(_06817_),
    .B(net275),
    .C(_06816_),
    .Y(_06819_));
 sky130_fd_sc_hd__o31a_1 _17364_ (.A1(net301),
    .A2(net300),
    .A3(_06805_),
    .B1(_06819_),
    .X(_06820_));
 sky130_fd_sc_hd__o22a_2 _17365_ (.A1(_05228_),
    .A2(_05230_),
    .B1(_06806_),
    .B2(_06818_),
    .X(_06821_));
 sky130_fd_sc_hd__or3_1 _17366_ (.A(net297),
    .B(_05232_),
    .C(_06820_),
    .X(_06822_));
 sky130_fd_sc_hd__a21o_1 _17367_ (.A1(_07044_),
    .A2(_06546_),
    .B1(_06547_),
    .X(_06823_));
 sky130_fd_sc_hd__o21a_1 _17368_ (.A1(_06229_),
    .A2(_06236_),
    .B1(_06548_),
    .X(_06824_));
 sky130_fd_sc_hd__a311oi_4 _17369_ (.A1(_06817_),
    .A2(net275),
    .A3(_06816_),
    .B1(_06806_),
    .C1(_07899_),
    .Y(_06825_));
 sky130_fd_sc_hd__o221ai_4 _17370_ (.A1(net369),
    .A2(_07866_),
    .B1(net275),
    .B2(_06805_),
    .C1(_06819_),
    .Y(_06827_));
 sky130_fd_sc_hd__a22oi_4 _17371_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_06807_),
    .B2(_06819_),
    .Y(_06828_));
 sky130_fd_sc_hd__o22ai_4 _17372_ (.A1(net390),
    .A2(net370),
    .B1(_06806_),
    .B2(_06818_),
    .Y(_06829_));
 sky130_fd_sc_hd__o21ai_2 _17373_ (.A1(_06549_),
    .A2(_06824_),
    .B1(_06827_),
    .Y(_06830_));
 sky130_fd_sc_hd__o211ai_4 _17374_ (.A1(_06549_),
    .A2(_06824_),
    .B1(_06827_),
    .C1(_06829_),
    .Y(_06831_));
 sky130_fd_sc_hd__o2bb2ai_4 _17375_ (.A1_N(_06548_),
    .A2_N(_06823_),
    .B1(_06825_),
    .B2(_06828_),
    .Y(_06832_));
 sky130_fd_sc_hd__o211ai_4 _17376_ (.A1(_06828_),
    .A2(_06830_),
    .B1(net274),
    .C1(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__o31a_2 _17377_ (.A1(net297),
    .A2(_05232_),
    .A3(_06820_),
    .B1(_06833_),
    .X(_06834_));
 sky130_fd_sc_hd__a31o_1 _17378_ (.A1(_06832_),
    .A2(net274),
    .A3(_06831_),
    .B1(_06821_),
    .X(_06835_));
 sky130_fd_sc_hd__a31o_1 _17379_ (.A1(_06832_),
    .A2(net274),
    .A3(_06831_),
    .B1(_07044_),
    .X(_06836_));
 sky130_fd_sc_hd__a311oi_4 _17380_ (.A1(_06832_),
    .A2(net274),
    .A3(_06831_),
    .B1(_06821_),
    .C1(_07044_),
    .Y(_06838_));
 sky130_fd_sc_hd__a22oi_4 _17381_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_06822_),
    .B2(_06833_),
    .Y(_06839_));
 sky130_fd_sc_hd__o21ai_1 _17382_ (.A1(_06945_),
    .A2(_06967_),
    .B1(_06835_),
    .Y(_06840_));
 sky130_fd_sc_hd__o211ai_2 _17383_ (.A1(_06836_),
    .A2(_06821_),
    .B1(_06620_),
    .C1(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__o21ai_1 _17384_ (.A1(_06838_),
    .A2(_06839_),
    .B1(_06619_),
    .Y(_06842_));
 sky130_fd_sc_hd__o211ai_4 _17385_ (.A1(_05481_),
    .A2(net269),
    .B1(_06841_),
    .C1(_06842_),
    .Y(_06843_));
 sky130_fd_sc_hd__a211o_1 _17386_ (.A1(_06822_),
    .A2(_06833_),
    .B1(_05481_),
    .C1(net269),
    .X(_06844_));
 sky130_fd_sc_hd__o31a_1 _17387_ (.A1(_05481_),
    .A2(net269),
    .A3(_06834_),
    .B1(_06843_),
    .X(_06845_));
 sky130_fd_sc_hd__o311a_1 _17388_ (.A1(_05481_),
    .A2(net269),
    .A3(_06834_),
    .B1(_06843_),
    .C1(_05754_),
    .X(_06846_));
 sky130_fd_sc_hd__a21oi_2 _17389_ (.A1(_06843_),
    .A2(_06844_),
    .B1(_06332_),
    .Y(_06847_));
 sky130_fd_sc_hd__a22o_1 _17390_ (.A1(_06256_),
    .A2(_06278_),
    .B1(_06843_),
    .B2(_06844_),
    .X(_06849_));
 sky130_fd_sc_hd__o221a_1 _17391_ (.A1(_06289_),
    .A2(_06310_),
    .B1(_05485_),
    .B2(_06834_),
    .C1(_06843_),
    .X(_06850_));
 sky130_fd_sc_hd__o221ai_4 _17392_ (.A1(_06289_),
    .A2(_06310_),
    .B1(_05485_),
    .B2(_06834_),
    .C1(_06843_),
    .Y(_06851_));
 sky130_fd_sc_hd__a22oi_2 _17393_ (.A1(_06559_),
    .A2(_06567_),
    .B1(_06573_),
    .B2(_05851_),
    .Y(_06852_));
 sky130_fd_sc_hd__a32o_1 _17394_ (.A1(_06571_),
    .A2(_05851_),
    .A3(_06264_),
    .B1(_06567_),
    .B2(_06559_),
    .X(_06853_));
 sky130_fd_sc_hd__o221ai_4 _17395_ (.A1(_05851_),
    .A2(_06573_),
    .B1(_06847_),
    .B2(_06850_),
    .C1(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__o21ai_4 _17396_ (.A1(_06575_),
    .A2(_06852_),
    .B1(_06851_),
    .Y(_06855_));
 sky130_fd_sc_hd__o211ai_1 _17397_ (.A1(_06575_),
    .A2(_06852_),
    .B1(_06851_),
    .C1(_06849_),
    .Y(_06856_));
 sky130_fd_sc_hd__a21oi_2 _17398_ (.A1(_06854_),
    .A2(_06856_),
    .B1(_05754_),
    .Y(_06857_));
 sky130_fd_sc_hd__o221ai_2 _17399_ (.A1(net266),
    .A2(_05751_),
    .B1(_06847_),
    .B2(_06855_),
    .C1(_06854_),
    .Y(_06858_));
 sky130_fd_sc_hd__o21ai_2 _17400_ (.A1(net241),
    .A2(_06845_),
    .B1(_06858_),
    .Y(_06860_));
 sky130_fd_sc_hd__nand4_2 _17401_ (.A(_06275_),
    .B(_06277_),
    .C(_06578_),
    .D(_06579_),
    .Y(_06861_));
 sky130_fd_sc_hd__o211ai_2 _17402_ (.A1(net387),
    .A2(_06581_),
    .B1(_06589_),
    .C1(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__o2111ai_4 _17403_ (.A1(net387),
    .A2(_06581_),
    .B1(_06589_),
    .C1(_05851_),
    .D1(_06861_),
    .Y(_06863_));
 sky130_fd_sc_hd__o21a_1 _17404_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_06862_),
    .X(_06864_));
 sky130_fd_sc_hd__o21ai_2 _17405_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_06862_),
    .Y(_06865_));
 sky130_fd_sc_hd__o211ai_2 _17406_ (.A1(net259),
    .A2(net256),
    .B1(_06863_),
    .C1(_06865_),
    .Y(_06866_));
 sky130_fd_sc_hd__and4_1 _17407_ (.A(_06860_),
    .B(_06863_),
    .C(_06865_),
    .D(_05996_),
    .X(_06867_));
 sky130_fd_sc_hd__nand4_2 _17408_ (.A(_06860_),
    .B(_06863_),
    .C(_06865_),
    .D(_05996_),
    .Y(_06868_));
 sky130_fd_sc_hd__o21ai_4 _17409_ (.A1(_06846_),
    .A2(_06857_),
    .B1(_06866_),
    .Y(_06869_));
 sky130_fd_sc_hd__inv_2 _17410_ (.A(_06869_),
    .Y(_06871_));
 sky130_fd_sc_hd__o31a_1 _17411_ (.A1(_06846_),
    .A2(_06857_),
    .A3(_06866_),
    .B1(_06869_),
    .X(_06872_));
 sky130_fd_sc_hd__nand2_1 _17412_ (.A(_06868_),
    .B(_06869_),
    .Y(_06873_));
 sky130_fd_sc_hd__nand2_1 _17413_ (.A(_06592_),
    .B(_06595_),
    .Y(_06874_));
 sky130_fd_sc_hd__o211ai_4 _17414_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_06592_),
    .C1(_06595_),
    .Y(_06875_));
 sky130_fd_sc_hd__o22ai_4 _17415_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_06591_),
    .B2(_06594_),
    .Y(_06876_));
 sky130_fd_sc_hd__nand3_1 _17416_ (.A(_06876_),
    .B(net212),
    .C(_06875_),
    .Y(_06877_));
 sky130_fd_sc_hd__a31o_1 _17417_ (.A1(_06876_),
    .A2(net212),
    .A3(_06875_),
    .B1(_06873_),
    .X(_06878_));
 sky130_fd_sc_hd__nand4_2 _17418_ (.A(_06873_),
    .B(_06875_),
    .C(_06876_),
    .D(net212),
    .Y(_06879_));
 sky130_fd_sc_hd__nand4_1 _17419_ (.A(net212),
    .B(_06872_),
    .C(_06875_),
    .D(_06876_),
    .Y(_06880_));
 sky130_fd_sc_hd__o21ai_1 _17420_ (.A1(_06867_),
    .A2(_06871_),
    .B1(_06877_),
    .Y(_06882_));
 sky130_fd_sc_hd__o211ai_2 _17421_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_06868_),
    .C1(_06869_),
    .Y(_06883_));
 sky130_fd_sc_hd__nand2_1 _17422_ (.A(_06880_),
    .B(_06882_),
    .Y(_06884_));
 sky130_fd_sc_hd__nand3_1 _17423_ (.A(_05250_),
    .B(_06878_),
    .C(_06879_),
    .Y(_06885_));
 sky130_fd_sc_hd__a21oi_2 _17424_ (.A1(_06878_),
    .A2(_06879_),
    .B1(_05250_),
    .Y(_06886_));
 sky130_fd_sc_hd__nand3_2 _17425_ (.A(_06882_),
    .B(net403),
    .C(_06880_),
    .Y(_06887_));
 sky130_fd_sc_hd__o31ai_2 _17426_ (.A1(_06601_),
    .A2(_03289_),
    .A3(_06600_),
    .B1(_06887_),
    .Y(_06888_));
 sky130_fd_sc_hd__a22o_1 _17427_ (.A1(net1),
    .A2(_06603_),
    .B1(_06885_),
    .B2(_06887_),
    .X(_06889_));
 sky130_fd_sc_hd__a31oi_1 _17428_ (.A1(_05250_),
    .A2(_06878_),
    .A3(_06879_),
    .B1(_06615_),
    .Y(_06890_));
 sky130_fd_sc_hd__a31o_1 _17429_ (.A1(_05250_),
    .A2(_06878_),
    .A3(_06879_),
    .B1(_06615_),
    .X(_06891_));
 sky130_fd_sc_hd__o211ai_2 _17430_ (.A1(_06886_),
    .A2(_06891_),
    .B1(_06612_),
    .C1(_06889_),
    .Y(_06893_));
 sky130_fd_sc_hd__or3_1 _17431_ (.A(_06608_),
    .B(net237),
    .C(_06884_),
    .X(_06894_));
 sky130_fd_sc_hd__o31a_1 _17432_ (.A1(_06608_),
    .A2(net237),
    .A3(_06884_),
    .B1(_06893_),
    .X(_06895_));
 sky130_fd_sc_hd__or4_4 _17433_ (.A(net40),
    .B(net41),
    .C(net42),
    .D(_05989_),
    .X(_06896_));
 sky130_fd_sc_hd__o311a_4 _17434_ (.A1(net41),
    .A2(net42),
    .A3(_06285_),
    .B1(net43),
    .C1(net409),
    .X(_06897_));
 sky130_fd_sc_hd__a21oi_4 _17435_ (.A1(_06896_),
    .A2(net409),
    .B1(net43),
    .Y(_06898_));
 sky130_fd_sc_hd__a21boi_4 _17436_ (.A1(_06896_),
    .A2(net409),
    .B1_N(net43),
    .Y(_06899_));
 sky130_fd_sc_hd__a21bo_4 _17437_ (.A1(_06896_),
    .A2(net409),
    .B1_N(net43),
    .X(_06900_));
 sky130_fd_sc_hd__and3b_4 _17438_ (.A_N(net43),
    .B(_06896_),
    .C(net409),
    .X(_06901_));
 sky130_fd_sc_hd__nand3b_4 _17439_ (.A_N(net43),
    .B(_06896_),
    .C(net409),
    .Y(_06902_));
 sky130_fd_sc_hd__nand2_8 _17440_ (.A(_06900_),
    .B(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__nor2_8 _17441_ (.A(net231),
    .B(net228),
    .Y(_06904_));
 sky130_fd_sc_hd__o2bb2a_1 _17442_ (.A1_N(_06893_),
    .A2_N(_06894_),
    .B1(_06904_),
    .B2(_03289_),
    .X(_06905_));
 sky130_fd_sc_hd__a21oi_1 _17443_ (.A1(_06893_),
    .A2(_06894_),
    .B1(_03289_),
    .Y(_06906_));
 sky130_fd_sc_hd__a31o_1 _17444_ (.A1(net1),
    .A2(_06895_),
    .A3(net208),
    .B1(_06905_),
    .X(_06907_));
 sky130_fd_sc_hd__xor2_1 _17445_ (.A(_06618_),
    .B(_06907_),
    .X(net75));
 sky130_fd_sc_hd__nor4_1 _17446_ (.A(_06003_),
    .B(_06299_),
    .C(_06616_),
    .D(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__a21oi_1 _17447_ (.A1(_07044_),
    .A2(_06835_),
    .B1(_06620_),
    .Y(_06909_));
 sky130_fd_sc_hd__o21ai_1 _17448_ (.A1(_06619_),
    .A2(_06838_),
    .B1(_06840_),
    .Y(_06910_));
 sky130_fd_sc_hd__o32ai_4 _17449_ (.A1(_06945_),
    .A2(_06967_),
    .A3(_06835_),
    .B1(_06620_),
    .B2(_06839_),
    .Y(_06911_));
 sky130_fd_sc_hd__or4_4 _17450_ (.A(net9),
    .B(net10),
    .C(net11),
    .D(_06008_),
    .X(_06913_));
 sky130_fd_sc_hd__and3b_4 _17451_ (.A_N(net13),
    .B(_06913_),
    .C(net410),
    .X(_06914_));
 sky130_fd_sc_hd__or3b_4 _17452_ (.A(_03399_),
    .B(net13),
    .C_N(_06913_),
    .X(_06915_));
 sky130_fd_sc_hd__a21boi_4 _17453_ (.A1(_06913_),
    .A2(net410),
    .B1_N(net13),
    .Y(_06916_));
 sky130_fd_sc_hd__a21bo_4 _17454_ (.A1(_06913_),
    .A2(net410),
    .B1_N(net13),
    .X(_06917_));
 sky130_fd_sc_hd__o311a_4 _17455_ (.A1(net10),
    .A2(net11),
    .A3(_06304_),
    .B1(net13),
    .C1(net410),
    .X(_06918_));
 sky130_fd_sc_hd__nand3_4 _17456_ (.A(_06913_),
    .B(net13),
    .C(net410),
    .Y(_06919_));
 sky130_fd_sc_hd__a21oi_4 _17457_ (.A1(_06913_),
    .A2(net410),
    .B1(net13),
    .Y(_06920_));
 sky130_fd_sc_hd__a21o_4 _17458_ (.A1(_06913_),
    .A2(net410),
    .B1(net13),
    .X(_06921_));
 sky130_fd_sc_hd__nand2_8 _17459_ (.A(_06919_),
    .B(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__nor2_8 _17460_ (.A(_06918_),
    .B(net249),
    .Y(_06924_));
 sky130_fd_sc_hd__or3_4 _17461_ (.A(_03178_),
    .B(_06918_),
    .C(_06920_),
    .X(_06925_));
 sky130_fd_sc_hd__o221a_1 _17462_ (.A1(_05130_),
    .A2(_05152_),
    .B1(_06914_),
    .B2(_06916_),
    .C1(net33),
    .X(_06926_));
 sky130_fd_sc_hd__and3_1 _17463_ (.A(net232),
    .B(net225),
    .C(net33),
    .X(_06927_));
 sky130_fd_sc_hd__or4_1 _17464_ (.A(_06918_),
    .B(_03178_),
    .C(net234),
    .D(_06920_),
    .X(_06928_));
 sky130_fd_sc_hd__o32a_2 _17465_ (.A1(_03178_),
    .A2(_06918_),
    .A3(_06920_),
    .B1(_06626_),
    .B2(_06627_),
    .X(_06929_));
 sky130_fd_sc_hd__a21oi_4 _17466_ (.A1(_06631_),
    .A2(net225),
    .B1(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__o211ai_4 _17467_ (.A1(_06327_),
    .A2(_06320_),
    .B1(_06324_),
    .C1(_06632_),
    .Y(_06931_));
 sky130_fd_sc_hd__o211ai_2 _17468_ (.A1(_06927_),
    .A2(_06929_),
    .B1(_06632_),
    .C1(_06635_),
    .Y(_06932_));
 sky130_fd_sc_hd__o211ai_4 _17469_ (.A1(net251),
    .A2(_06631_),
    .B1(_06930_),
    .C1(_06931_),
    .Y(_06933_));
 sky130_fd_sc_hd__o32a_2 _17470_ (.A1(_03178_),
    .A2(_06918_),
    .A3(_06920_),
    .B1(_05130_),
    .B2(_05152_),
    .X(_06935_));
 sky130_fd_sc_hd__a31o_1 _17471_ (.A1(_06921_),
    .A2(net33),
    .A3(_06919_),
    .B1(net405),
    .X(_06936_));
 sky130_fd_sc_hd__a21oi_1 _17472_ (.A1(_06932_),
    .A2(_06933_),
    .B1(_05185_),
    .Y(_06937_));
 sky130_fd_sc_hd__a21o_1 _17473_ (.A1(_06932_),
    .A2(_06933_),
    .B1(_05185_),
    .X(_06938_));
 sky130_fd_sc_hd__a21o_1 _17474_ (.A1(_05185_),
    .A2(_06925_),
    .B1(_06937_),
    .X(_06939_));
 sky130_fd_sc_hd__a31oi_4 _17475_ (.A1(_06647_),
    .A2(_06648_),
    .A3(_06340_),
    .B1(_06645_),
    .Y(_06940_));
 sky130_fd_sc_hd__a311oi_2 _17476_ (.A1(_06932_),
    .A2(_06933_),
    .A3(net405),
    .B1(net251),
    .C1(_06926_),
    .Y(_06941_));
 sky130_fd_sc_hd__a311o_2 _17477_ (.A1(_06932_),
    .A2(_06933_),
    .A3(net405),
    .B1(net251),
    .C1(_06926_),
    .X(_06942_));
 sky130_fd_sc_hd__o21ai_2 _17478_ (.A1(_06305_),
    .A2(net283),
    .B1(_06938_),
    .Y(_06943_));
 sky130_fd_sc_hd__nor3_1 _17479_ (.A(_06314_),
    .B(_06935_),
    .C(_06937_),
    .Y(_06944_));
 sky130_fd_sc_hd__a211o_1 _17480_ (.A1(_06306_),
    .A2(_06308_),
    .B1(_06935_),
    .C1(_06937_),
    .X(_06946_));
 sky130_fd_sc_hd__o21ai_4 _17481_ (.A1(_06935_),
    .A2(_06943_),
    .B1(_06942_),
    .Y(_06947_));
 sky130_fd_sc_hd__o221ai_2 _17482_ (.A1(net254),
    .A2(_06641_),
    .B1(_06941_),
    .B2(_06944_),
    .C1(_06649_),
    .Y(_06948_));
 sky130_fd_sc_hd__a21oi_4 _17483_ (.A1(_06646_),
    .A2(_06649_),
    .B1(_06947_),
    .Y(_06949_));
 sky130_fd_sc_hd__and3_1 _17484_ (.A(_06938_),
    .B(_05392_),
    .C(_06936_),
    .X(_06950_));
 sky130_fd_sc_hd__o21ai_2 _17485_ (.A1(net402),
    .A2(_05370_),
    .B1(_06948_),
    .Y(_06951_));
 sky130_fd_sc_hd__o22ai_2 _17486_ (.A1(net388),
    .A2(_06939_),
    .B1(_06949_),
    .B2(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__o22a_2 _17487_ (.A1(net388),
    .A2(_06939_),
    .B1(_06949_),
    .B2(_06951_),
    .X(_06953_));
 sky130_fd_sc_hd__and3_2 _17488_ (.A(_06952_),
    .B(_05709_),
    .C(_05687_),
    .X(_06954_));
 sky130_fd_sc_hd__o21ai_4 _17489_ (.A1(_06009_),
    .A2(_06010_),
    .B1(_06952_),
    .Y(_06955_));
 sky130_fd_sc_hd__inv_2 _17490_ (.A(_06955_),
    .Y(_06957_));
 sky130_fd_sc_hd__o21ai_2 _17491_ (.A1(_06949_),
    .A2(_06951_),
    .B1(net254),
    .Y(_06958_));
 sky130_fd_sc_hd__o21ai_4 _17492_ (.A1(_06950_),
    .A2(_06958_),
    .B1(_06955_),
    .Y(_06959_));
 sky130_fd_sc_hd__a31oi_4 _17493_ (.A1(_06660_),
    .A2(_06668_),
    .A3(_06670_),
    .B1(_06657_),
    .Y(_06960_));
 sky130_fd_sc_hd__o311a_4 _17494_ (.A1(_05765_),
    .A2(net289),
    .A3(_06654_),
    .B1(_06674_),
    .C1(_06959_),
    .X(_06961_));
 sky130_fd_sc_hd__o21ai_4 _17495_ (.A1(_06959_),
    .A2(_06960_),
    .B1(net359),
    .Y(_06962_));
 sky130_fd_sc_hd__o22ai_4 _17496_ (.A1(net359),
    .A2(_06953_),
    .B1(_06961_),
    .B2(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__and3_1 _17497_ (.A(_06804_),
    .B(_06826_),
    .C(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__or3b_2 _17498_ (.A(net379),
    .B(net378),
    .C_N(_06963_),
    .X(_06965_));
 sky130_fd_sc_hd__o21a_1 _17499_ (.A1(_05760_),
    .A2(net290),
    .B1(_06963_),
    .X(_06966_));
 sky130_fd_sc_hd__o21ai_4 _17500_ (.A1(_05760_),
    .A2(net290),
    .B1(_06963_),
    .Y(_06968_));
 sky130_fd_sc_hd__o21ai_4 _17501_ (.A1(_06961_),
    .A2(_06962_),
    .B1(net262),
    .Y(_06969_));
 sky130_fd_sc_hd__o221a_1 _17502_ (.A1(net359),
    .A2(_06953_),
    .B1(_06961_),
    .B2(_06962_),
    .C1(net262),
    .X(_06970_));
 sky130_fd_sc_hd__o221ai_4 _17503_ (.A1(net359),
    .A2(_06953_),
    .B1(_06961_),
    .B2(_06962_),
    .C1(net262),
    .Y(_06971_));
 sky130_fd_sc_hd__o21a_1 _17504_ (.A1(_06954_),
    .A2(_06969_),
    .B1(_06968_),
    .X(_06972_));
 sky130_fd_sc_hd__o21ai_4 _17505_ (.A1(_06954_),
    .A2(_06969_),
    .B1(_06968_),
    .Y(_06973_));
 sky130_fd_sc_hd__o211a_1 _17506_ (.A1(_06071_),
    .A2(_06080_),
    .B1(_06078_),
    .C1(_05831_),
    .X(_06974_));
 sky130_fd_sc_hd__o2111ai_1 _17507_ (.A1(_06071_),
    .A2(_06080_),
    .B1(_06078_),
    .C1(_05813_),
    .D1(_05815_),
    .Y(_06975_));
 sky130_fd_sc_hd__nor3_2 _17508_ (.A(_06381_),
    .B(_06383_),
    .C(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__nand4b_2 _17509_ (.A_N(_05827_),
    .B(_06382_),
    .C(_06974_),
    .D(_06384_),
    .Y(_06977_));
 sky130_fd_sc_hd__nand2_1 _17510_ (.A(_06976_),
    .B(_06685_),
    .Y(_06979_));
 sky130_fd_sc_hd__nand3_2 _17511_ (.A(_06685_),
    .B(_06687_),
    .C(_06976_),
    .Y(_06980_));
 sky130_fd_sc_hd__nor3_2 _17512_ (.A(_06977_),
    .B(_06686_),
    .C(_06684_),
    .Y(_06981_));
 sky130_fd_sc_hd__nand3b_1 _17513_ (.A_N(_06977_),
    .B(_06687_),
    .C(_06685_),
    .Y(_06982_));
 sky130_fd_sc_hd__a21oi_2 _17514_ (.A1(_06976_),
    .A2(_06685_),
    .B1(_06686_),
    .Y(_06983_));
 sky130_fd_sc_hd__o211a_1 _17515_ (.A1(_06684_),
    .A2(_06682_),
    .B1(_06979_),
    .C1(_06687_),
    .X(_06984_));
 sky130_fd_sc_hd__o211ai_4 _17516_ (.A1(_06684_),
    .A2(_06682_),
    .B1(_06979_),
    .C1(_06687_),
    .Y(_06985_));
 sky130_fd_sc_hd__a21oi_2 _17517_ (.A1(_06688_),
    .A2(_06983_),
    .B1(_06981_),
    .Y(_06986_));
 sky130_fd_sc_hd__o2bb2ai_4 _17518_ (.A1_N(_06983_),
    .A2_N(_06688_),
    .B1(_05827_),
    .B2(_06980_),
    .Y(_06987_));
 sky130_fd_sc_hd__o211ai_4 _17519_ (.A1(_05827_),
    .A2(_06980_),
    .B1(_06985_),
    .C1(_06973_),
    .Y(_06988_));
 sky130_fd_sc_hd__nand2_1 _17520_ (.A(_06987_),
    .B(_06972_),
    .Y(_06990_));
 sky130_fd_sc_hd__a211oi_2 _17521_ (.A1(_06688_),
    .A2(_06983_),
    .B1(_06981_),
    .C1(_06973_),
    .Y(_06991_));
 sky130_fd_sc_hd__nand4_1 _17522_ (.A(_06968_),
    .B(_06971_),
    .C(_06982_),
    .D(_06985_),
    .Y(_06992_));
 sky130_fd_sc_hd__o22ai_1 _17523_ (.A1(_06966_),
    .A2(_06970_),
    .B1(_06981_),
    .B2(_06984_),
    .Y(_06993_));
 sky130_fd_sc_hd__o22ai_2 _17524_ (.A1(net379),
    .A2(net378),
    .B1(_06972_),
    .B2(_06986_),
    .Y(_06994_));
 sky130_fd_sc_hd__nand3_1 _17525_ (.A(_06993_),
    .B(net357),
    .C(_06992_),
    .Y(_06995_));
 sky130_fd_sc_hd__o221a_1 _17526_ (.A1(net359),
    .A2(_06953_),
    .B1(_06961_),
    .B2(_06962_),
    .C1(_06848_),
    .X(_06996_));
 sky130_fd_sc_hd__nand3_1 _17527_ (.A(_06990_),
    .B(net357),
    .C(_06988_),
    .Y(_06997_));
 sky130_fd_sc_hd__a31o_1 _17528_ (.A1(_06990_),
    .A2(net357),
    .A3(_06988_),
    .B1(_06996_),
    .X(_06998_));
 sky130_fd_sc_hd__inv_2 _17529_ (.A(_06998_),
    .Y(_06999_));
 sky130_fd_sc_hd__o211a_2 _17530_ (.A1(_06963_),
    .A2(net357),
    .B1(_07724_),
    .C1(_06997_),
    .X(_07001_));
 sky130_fd_sc_hd__a311o_2 _17531_ (.A1(_06990_),
    .A2(net357),
    .A3(_06988_),
    .B1(_06996_),
    .C1(net356),
    .X(_07002_));
 sky130_fd_sc_hd__a31oi_1 _17532_ (.A1(_06993_),
    .A2(net357),
    .A3(_06992_),
    .B1(net291),
    .Y(_07003_));
 sky130_fd_sc_hd__o22ai_4 _17533_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_06991_),
    .B2(_06994_),
    .Y(_07004_));
 sky130_fd_sc_hd__o211ai_4 _17534_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_06965_),
    .C1(_06995_),
    .Y(_07005_));
 sky130_fd_sc_hd__a311oi_2 _17535_ (.A1(_06990_),
    .A2(net357),
    .A3(_06988_),
    .B1(_06996_),
    .C1(net267),
    .Y(_07006_));
 sky130_fd_sc_hd__o211ai_4 _17536_ (.A1(_06963_),
    .A2(net357),
    .B1(net291),
    .C1(_06997_),
    .Y(_07007_));
 sky130_fd_sc_hd__a21oi_1 _17537_ (.A1(net293),
    .A2(_06691_),
    .B1(_06695_),
    .Y(_07008_));
 sky130_fd_sc_hd__a21o_1 _17538_ (.A1(_06695_),
    .A2(_06697_),
    .B1(_06698_),
    .X(_07009_));
 sky130_fd_sc_hd__a21oi_1 _17539_ (.A1(_06695_),
    .A2(_06697_),
    .B1(_06698_),
    .Y(_07010_));
 sky130_fd_sc_hd__a21oi_1 _17540_ (.A1(_07005_),
    .A2(_07007_),
    .B1(_07009_),
    .Y(_07012_));
 sky130_fd_sc_hd__o2bb2ai_2 _17541_ (.A1_N(_07005_),
    .A2_N(_07007_),
    .B1(_07008_),
    .B2(_06696_),
    .Y(_07013_));
 sky130_fd_sc_hd__o211a_1 _17542_ (.A1(_06964_),
    .A2(_07004_),
    .B1(_07007_),
    .C1(_07009_),
    .X(_07014_));
 sky130_fd_sc_hd__nand3_2 _17543_ (.A(_07005_),
    .B(_07007_),
    .C(_07009_),
    .Y(_07015_));
 sky130_fd_sc_hd__nand3_2 _17544_ (.A(_07013_),
    .B(_07015_),
    .C(net355),
    .Y(_07016_));
 sky130_fd_sc_hd__o22ai_4 _17545_ (.A1(net373),
    .A2(net371),
    .B1(_07012_),
    .B2(_07014_),
    .Y(_07017_));
 sky130_fd_sc_hd__a31o_2 _17546_ (.A1(_07013_),
    .A2(_07015_),
    .A3(net355),
    .B1(_07001_),
    .X(_07018_));
 sky130_fd_sc_hd__a2bb2oi_4 _17547_ (.A1_N(_05242_),
    .A2_N(net314),
    .B1(_07002_),
    .B2(_07016_),
    .Y(_07019_));
 sky130_fd_sc_hd__o221ai_4 _17548_ (.A1(_05242_),
    .A2(net314),
    .B1(_06999_),
    .B2(net355),
    .C1(_07017_),
    .Y(_07020_));
 sky130_fd_sc_hd__a31oi_1 _17549_ (.A1(_07013_),
    .A2(_07015_),
    .A3(net355),
    .B1(net293),
    .Y(_07021_));
 sky130_fd_sc_hd__a31o_2 _17550_ (.A1(_07013_),
    .A2(_07015_),
    .A3(net355),
    .B1(net293),
    .X(_07023_));
 sky130_fd_sc_hd__o211a_1 _17551_ (.A1(net355),
    .A2(_06998_),
    .B1(net295),
    .C1(_07016_),
    .X(_07024_));
 sky130_fd_sc_hd__a311o_1 _17552_ (.A1(_07013_),
    .A2(_07015_),
    .A3(net355),
    .B1(net293),
    .C1(_07001_),
    .X(_07025_));
 sky130_fd_sc_hd__a21oi_1 _17553_ (.A1(_07002_),
    .A2(_07021_),
    .B1(_07019_),
    .Y(_07026_));
 sky130_fd_sc_hd__o32a_1 _17554_ (.A1(_04206_),
    .A2(_04216_),
    .A3(_06708_),
    .B1(_06712_),
    .B2(_06713_),
    .X(_07027_));
 sky130_fd_sc_hd__o22ai_4 _17555_ (.A1(net299),
    .A2(_06708_),
    .B1(_06712_),
    .B2(_06713_),
    .Y(_07028_));
 sky130_fd_sc_hd__a21oi_1 _17556_ (.A1(_07020_),
    .A2(_07025_),
    .B1(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__o21ai_4 _17557_ (.A1(_07019_),
    .A2(_07024_),
    .B1(_07027_),
    .Y(_07030_));
 sky130_fd_sc_hd__o211a_1 _17558_ (.A1(_07001_),
    .A2(_07023_),
    .B1(_07028_),
    .C1(_07020_),
    .X(_07031_));
 sky130_fd_sc_hd__o211ai_4 _17559_ (.A1(_07001_),
    .A2(_07023_),
    .B1(_07028_),
    .C1(_07020_),
    .Y(_07032_));
 sky130_fd_sc_hd__o22ai_2 _17560_ (.A1(net353),
    .A2(net352),
    .B1(_07029_),
    .B2(_07031_),
    .Y(_07034_));
 sky130_fd_sc_hd__o311a_2 _17561_ (.A1(net373),
    .A2(_06999_),
    .A3(net371),
    .B1(_08732_),
    .C1(_07017_),
    .X(_07035_));
 sky130_fd_sc_hd__a211o_1 _17562_ (.A1(_07002_),
    .A2(_07016_),
    .B1(net353),
    .C1(net352),
    .X(_07036_));
 sky130_fd_sc_hd__nand3_2 _17563_ (.A(_07030_),
    .B(_07032_),
    .C(net338),
    .Y(_07037_));
 sky130_fd_sc_hd__a31o_1 _17564_ (.A1(_07030_),
    .A2(_07032_),
    .A3(net338),
    .B1(_07035_),
    .X(_07038_));
 sky130_fd_sc_hd__a31oi_4 _17565_ (.A1(_07030_),
    .A2(_07032_),
    .A3(net338),
    .B1(_07035_),
    .Y(_07039_));
 sky130_fd_sc_hd__a2bb2oi_2 _17566_ (.A1_N(net339),
    .A2_N(_04184_),
    .B1(_07036_),
    .B2(_07037_),
    .Y(_07040_));
 sky130_fd_sc_hd__o221ai_4 _17567_ (.A1(net339),
    .A2(_04184_),
    .B1(_07018_),
    .B2(net338),
    .C1(_07034_),
    .Y(_07041_));
 sky130_fd_sc_hd__a311oi_4 _17568_ (.A1(_07030_),
    .A2(_07032_),
    .A3(net338),
    .B1(_07035_),
    .C1(net298),
    .Y(_07042_));
 sky130_fd_sc_hd__o211ai_4 _17569_ (.A1(_04206_),
    .A2(_04216_),
    .B1(_07036_),
    .C1(_07037_),
    .Y(_07043_));
 sky130_fd_sc_hd__o22a_1 _17570_ (.A1(_06717_),
    .A2(_06728_),
    .B1(_06725_),
    .B2(_06724_),
    .X(_07045_));
 sky130_fd_sc_hd__o22ai_4 _17571_ (.A1(_06717_),
    .A2(_06728_),
    .B1(_06725_),
    .B2(_06724_),
    .Y(_07046_));
 sky130_fd_sc_hd__nand3_1 _17572_ (.A(_07041_),
    .B(_07043_),
    .C(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__o21ai_1 _17573_ (.A1(_07040_),
    .A2(_07042_),
    .B1(_07045_),
    .Y(_07048_));
 sky130_fd_sc_hd__o211ai_4 _17574_ (.A1(_09785_),
    .A2(net349),
    .B1(_07047_),
    .C1(_07048_),
    .Y(_07049_));
 sky130_fd_sc_hd__o221a_2 _17575_ (.A1(_09763_),
    .A2(_09774_),
    .B1(_07018_),
    .B2(net338),
    .C1(_07034_),
    .X(_07050_));
 sky130_fd_sc_hd__or3_1 _17576_ (.A(net350),
    .B(net349),
    .C(_07039_),
    .X(_07051_));
 sky130_fd_sc_hd__o21ai_4 _17577_ (.A1(_07040_),
    .A2(_07042_),
    .B1(_07046_),
    .Y(_07052_));
 sky130_fd_sc_hd__nand3_4 _17578_ (.A(_07041_),
    .B(_07045_),
    .C(_07043_),
    .Y(_07053_));
 sky130_fd_sc_hd__nand3_2 _17579_ (.A(_07052_),
    .B(_07053_),
    .C(net337),
    .Y(_07054_));
 sky130_fd_sc_hd__o31a_2 _17580_ (.A1(net350),
    .A2(net349),
    .A3(_07039_),
    .B1(_07054_),
    .X(_07056_));
 sky130_fd_sc_hd__a311o_1 _17581_ (.A1(_07052_),
    .A2(_07053_),
    .A3(net336),
    .B1(net334),
    .C1(_07050_),
    .X(_07057_));
 sky130_fd_sc_hd__a22oi_4 _17582_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_07051_),
    .B2(_07054_),
    .Y(_07058_));
 sky130_fd_sc_hd__o2111ai_4 _17583_ (.A1(net337),
    .A2(_07038_),
    .B1(_07049_),
    .C1(_02104_),
    .D1(_02126_),
    .Y(_07059_));
 sky130_fd_sc_hd__a31o_1 _17584_ (.A1(_07052_),
    .A2(_07053_),
    .A3(net337),
    .B1(_02148_),
    .X(_07060_));
 sky130_fd_sc_hd__a311oi_4 _17585_ (.A1(_07052_),
    .A2(_07053_),
    .A3(net336),
    .B1(_02148_),
    .C1(_07050_),
    .Y(_07061_));
 sky130_fd_sc_hd__o211ai_4 _17586_ (.A1(net337),
    .A2(_07039_),
    .B1(_02137_),
    .C1(_07054_),
    .Y(_07062_));
 sky130_fd_sc_hd__nand4_2 _17587_ (.A(_05889_),
    .B(_05893_),
    .C(_06151_),
    .D(_06153_),
    .Y(_07063_));
 sky130_fd_sc_hd__a21oi_2 _17588_ (.A1(net325),
    .A2(_06457_),
    .B1(_07063_),
    .Y(_07064_));
 sky130_fd_sc_hd__nor3_1 _17589_ (.A(_06461_),
    .B(_07063_),
    .C(_06463_),
    .Y(_07065_));
 sky130_fd_sc_hd__nand3_1 _17590_ (.A(_07064_),
    .B(_06743_),
    .C(_06462_),
    .Y(_07067_));
 sky130_fd_sc_hd__o211a_1 _17591_ (.A1(_06748_),
    .A2(_06742_),
    .B1(_06745_),
    .C1(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__o211ai_4 _17592_ (.A1(_06748_),
    .A2(_06742_),
    .B1(_06745_),
    .C1(_07067_),
    .Y(_07069_));
 sky130_fd_sc_hd__nand4_4 _17593_ (.A(_06462_),
    .B(_07064_),
    .C(_06743_),
    .D(_05890_),
    .Y(_07070_));
 sky130_fd_sc_hd__nand4_4 _17594_ (.A(_06743_),
    .B(_07065_),
    .C(_06745_),
    .D(_05890_),
    .Y(_07071_));
 sky130_fd_sc_hd__o21ai_4 _17595_ (.A1(_06744_),
    .A2(_07070_),
    .B1(_07069_),
    .Y(_07072_));
 sky130_fd_sc_hd__o211ai_1 _17596_ (.A1(_07060_),
    .A2(_07050_),
    .B1(_07059_),
    .C1(_07072_),
    .Y(_07073_));
 sky130_fd_sc_hd__o221ai_1 _17597_ (.A1(_06744_),
    .A2(_07070_),
    .B1(_07061_),
    .B2(_07058_),
    .C1(_07069_),
    .Y(_07074_));
 sky130_fd_sc_hd__nand3_1 _17598_ (.A(_07073_),
    .B(_07074_),
    .C(net334),
    .Y(_07075_));
 sky130_fd_sc_hd__o211a_1 _17599_ (.A1(net337),
    .A2(_07038_),
    .B1(_07049_),
    .C1(_11079_),
    .X(_07076_));
 sky130_fd_sc_hd__or3_1 _17600_ (.A(net347),
    .B(net346),
    .C(_07056_),
    .X(_07078_));
 sky130_fd_sc_hd__o21ai_1 _17601_ (.A1(_06744_),
    .A2(_07070_),
    .B1(_07062_),
    .Y(_07079_));
 sky130_fd_sc_hd__o211ai_4 _17602_ (.A1(_07070_),
    .A2(_06744_),
    .B1(_07062_),
    .C1(_07069_),
    .Y(_07080_));
 sky130_fd_sc_hd__nand4_4 _17603_ (.A(_07059_),
    .B(_07062_),
    .C(_07069_),
    .D(_07071_),
    .Y(_07081_));
 sky130_fd_sc_hd__o21ai_4 _17604_ (.A1(_07058_),
    .A2(_07061_),
    .B1(_07072_),
    .Y(_07082_));
 sky130_fd_sc_hd__nand3_2 _17605_ (.A(_07082_),
    .B(net334),
    .C(_07081_),
    .Y(_07083_));
 sky130_fd_sc_hd__a31oi_4 _17606_ (.A1(_07082_),
    .A2(net334),
    .A3(_07081_),
    .B1(_07076_),
    .Y(_07084_));
 sky130_fd_sc_hd__and3_2 _17607_ (.A(_12703_),
    .B(_07057_),
    .C(_07075_),
    .X(_07085_));
 sky130_fd_sc_hd__or3_1 _17608_ (.A(_12670_),
    .B(_12681_),
    .C(_07084_),
    .X(_07086_));
 sky130_fd_sc_hd__a31oi_2 _17609_ (.A1(_07082_),
    .A2(net334),
    .A3(_07081_),
    .B1(net319),
    .Y(_07087_));
 sky130_fd_sc_hd__o211a_2 _17610_ (.A1(net334),
    .A2(_07056_),
    .B1(net320),
    .C1(_07083_),
    .X(_07089_));
 sky130_fd_sc_hd__o211ai_4 _17611_ (.A1(net334),
    .A2(_07056_),
    .B1(net320),
    .C1(_07083_),
    .Y(_07090_));
 sky130_fd_sc_hd__o211ai_4 _17612_ (.A1(_00174_),
    .A2(_00196_),
    .B1(_07057_),
    .C1(_07075_),
    .Y(_07091_));
 sky130_fd_sc_hd__o211a_1 _17613_ (.A1(_12888_),
    .A2(_06753_),
    .B1(_06490_),
    .C1(_06477_),
    .X(_07092_));
 sky130_fd_sc_hd__a21oi_2 _17614_ (.A1(_06477_),
    .A2(_06490_),
    .B1(_06757_),
    .Y(_07093_));
 sky130_fd_sc_hd__o31ai_2 _17615_ (.A1(_06476_),
    .A2(_06756_),
    .A3(_06759_),
    .B1(_06758_),
    .Y(_07094_));
 sky130_fd_sc_hd__a21boi_1 _17616_ (.A1(_07090_),
    .A2(_07091_),
    .B1_N(_07094_),
    .Y(_07095_));
 sky130_fd_sc_hd__o2bb2ai_4 _17617_ (.A1_N(_07090_),
    .A2_N(_07091_),
    .B1(_07092_),
    .B2(_06757_),
    .Y(_07096_));
 sky130_fd_sc_hd__o22ai_1 _17618_ (.A1(_06759_),
    .A2(_07093_),
    .B1(net320),
    .B2(_07084_),
    .Y(_07097_));
 sky130_fd_sc_hd__o211ai_4 _17619_ (.A1(_06759_),
    .A2(_07093_),
    .B1(_07091_),
    .C1(_07090_),
    .Y(_07098_));
 sky130_fd_sc_hd__o22ai_2 _17620_ (.A1(_12670_),
    .A2(_12681_),
    .B1(_07089_),
    .B2(_07097_),
    .Y(_07100_));
 sky130_fd_sc_hd__nand3_2 _17621_ (.A(_07096_),
    .B(_07098_),
    .C(net312),
    .Y(_07101_));
 sky130_fd_sc_hd__a31oi_4 _17622_ (.A1(_07096_),
    .A2(_07098_),
    .A3(net312),
    .B1(_07085_),
    .Y(_07102_));
 sky130_fd_sc_hd__o22ai_4 _17623_ (.A1(net312),
    .A2(_07084_),
    .B1(_07095_),
    .B2(_07100_),
    .Y(_07103_));
 sky130_fd_sc_hd__o221a_1 _17624_ (.A1(_06498_),
    .A2(_06501_),
    .B1(net331),
    .B2(_06770_),
    .C1(_06496_),
    .X(_07104_));
 sky130_fd_sc_hd__o311a_1 _17625_ (.A1(_06189_),
    .A2(_06495_),
    .A3(_06500_),
    .B1(_06774_),
    .C1(_06499_),
    .X(_07105_));
 sky130_fd_sc_hd__o21ai_2 _17626_ (.A1(_06779_),
    .A2(_06773_),
    .B1(_06776_),
    .Y(_07106_));
 sky130_fd_sc_hd__a311oi_4 _17627_ (.A1(_07096_),
    .A2(_07098_),
    .A3(net312),
    .B1(net325),
    .C1(_07085_),
    .Y(_07107_));
 sky130_fd_sc_hd__o221ai_4 _17628_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_07084_),
    .B2(net312),
    .C1(_07101_),
    .Y(_07108_));
 sky130_fd_sc_hd__a2bb2oi_4 _17629_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_07086_),
    .B2(_07101_),
    .Y(_07109_));
 sky130_fd_sc_hd__o21ai_2 _17630_ (.A1(_12845_),
    .A2(_12856_),
    .B1(_07103_),
    .Y(_07111_));
 sky130_fd_sc_hd__o2111ai_1 _17631_ (.A1(_06779_),
    .A2(_06773_),
    .B1(_06776_),
    .C1(_07108_),
    .D1(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__o22ai_1 _17632_ (.A1(_06775_),
    .A2(_07105_),
    .B1(_07107_),
    .B2(_07109_),
    .Y(_07113_));
 sky130_fd_sc_hd__nand3_1 _17633_ (.A(_07112_),
    .B(_07113_),
    .C(net309),
    .Y(_07114_));
 sky130_fd_sc_hd__and3_1 _17634_ (.A(_00022_),
    .B(_00044_),
    .C(_07103_),
    .X(_07115_));
 sky130_fd_sc_hd__o21ai_1 _17635_ (.A1(_12888_),
    .A2(_07102_),
    .B1(_07106_),
    .Y(_07116_));
 sky130_fd_sc_hd__o211ai_4 _17636_ (.A1(_06775_),
    .A2(_07105_),
    .B1(_07108_),
    .C1(_07111_),
    .Y(_07117_));
 sky130_fd_sc_hd__o22ai_4 _17637_ (.A1(_06773_),
    .A2(_07104_),
    .B1(_07107_),
    .B2(_07109_),
    .Y(_07118_));
 sky130_fd_sc_hd__o221ai_4 _17638_ (.A1(net324),
    .A2(_00033_),
    .B1(_07107_),
    .B2(_07116_),
    .C1(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__a31o_1 _17639_ (.A1(_07117_),
    .A2(_07118_),
    .A3(net310),
    .B1(_07115_),
    .X(_07120_));
 sky130_fd_sc_hd__a31oi_4 _17640_ (.A1(_07117_),
    .A2(_07118_),
    .A3(net310),
    .B1(_07115_),
    .Y(_07122_));
 sky130_fd_sc_hd__o211ai_4 _17641_ (.A1(_07103_),
    .A2(net309),
    .B1(net330),
    .C1(_07114_),
    .Y(_07123_));
 sky130_fd_sc_hd__o211a_1 _17642_ (.A1(net309),
    .A2(_07102_),
    .B1(net331),
    .C1(_07119_),
    .X(_07124_));
 sky130_fd_sc_hd__o211ai_4 _17643_ (.A1(net309),
    .A2(_07102_),
    .B1(net331),
    .C1(_07119_),
    .Y(_07125_));
 sky130_fd_sc_hd__o311a_1 _17644_ (.A1(_06201_),
    .A2(_06514_),
    .A3(_06518_),
    .B1(_06790_),
    .C1(_06517_),
    .X(_07126_));
 sky130_fd_sc_hd__o21ai_2 _17645_ (.A1(_06791_),
    .A2(_06794_),
    .B1(_06790_),
    .Y(_07127_));
 sky130_fd_sc_hd__o2bb2ai_2 _17646_ (.A1_N(_07123_),
    .A2_N(_07125_),
    .B1(_07126_),
    .B2(_06791_),
    .Y(_07128_));
 sky130_fd_sc_hd__nand3_2 _17647_ (.A(_07123_),
    .B(_07125_),
    .C(_07127_),
    .Y(_07129_));
 sky130_fd_sc_hd__a31oi_2 _17648_ (.A1(_07123_),
    .A2(_07125_),
    .A3(_07127_),
    .B1(_01973_),
    .Y(_07130_));
 sky130_fd_sc_hd__nand3_4 _17649_ (.A(_07128_),
    .B(_07129_),
    .C(_01962_),
    .Y(_07131_));
 sky130_fd_sc_hd__or3_1 _17650_ (.A(net305),
    .B(net303),
    .C(_07122_),
    .X(_07133_));
 sky130_fd_sc_hd__o2bb2ai_4 _17651_ (.A1_N(_07130_),
    .A2_N(_07128_),
    .B1(_07122_),
    .B2(_01962_),
    .Y(_07134_));
 sky130_fd_sc_hd__a22oi_2 _17652_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_07131_),
    .B2(_07133_),
    .Y(_07135_));
 sky130_fd_sc_hd__a22o_2 _17653_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_07131_),
    .B2(_07133_),
    .X(_07136_));
 sky130_fd_sc_hd__o221a_2 _17654_ (.A1(_09971_),
    .A2(_09993_),
    .B1(net280),
    .B2(_07122_),
    .C1(_07131_),
    .X(_07137_));
 sky130_fd_sc_hd__o221ai_4 _17655_ (.A1(_09971_),
    .A2(_09993_),
    .B1(net280),
    .B2(_07122_),
    .C1(_07131_),
    .Y(_07138_));
 sky130_fd_sc_hd__o32a_2 _17656_ (.A1(_08863_),
    .A2(_06805_),
    .A3(net366),
    .B1(_06809_),
    .B2(_06808_),
    .X(_07139_));
 sky130_fd_sc_hd__o21ai_2 _17657_ (.A1(_06808_),
    .A2(_06809_),
    .B1(_06812_),
    .Y(_07140_));
 sky130_fd_sc_hd__o21ai_1 _17658_ (.A1(_07135_),
    .A2(_07137_),
    .B1(_07139_),
    .Y(_07141_));
 sky130_fd_sc_hd__nand3_1 _17659_ (.A(_07136_),
    .B(_07138_),
    .C(_07140_),
    .Y(_07142_));
 sky130_fd_sc_hd__nand3_1 _17660_ (.A(_07136_),
    .B(_07138_),
    .C(_07139_),
    .Y(_07144_));
 sky130_fd_sc_hd__o21ai_1 _17661_ (.A1(_07135_),
    .A2(_07137_),
    .B1(_07140_),
    .Y(_07145_));
 sky130_fd_sc_hd__o211ai_4 _17662_ (.A1(net301),
    .A2(net300),
    .B1(_07144_),
    .C1(_07145_),
    .Y(_07146_));
 sky130_fd_sc_hd__a211o_1 _17663_ (.A1(_07131_),
    .A2(_07133_),
    .B1(net301),
    .C1(net300),
    .X(_07147_));
 sky130_fd_sc_hd__nand3_2 _17664_ (.A(_07141_),
    .B(_07142_),
    .C(net275),
    .Y(_07148_));
 sky130_fd_sc_hd__o311a_2 _17665_ (.A1(net301),
    .A2(_07134_),
    .A3(net300),
    .B1(_05234_),
    .C1(_07146_),
    .X(_07149_));
 sky130_fd_sc_hd__a211o_1 _17666_ (.A1(_07147_),
    .A2(_07148_),
    .B1(net297),
    .C1(_05232_),
    .X(_07150_));
 sky130_fd_sc_hd__nand3_2 _17667_ (.A(_07148_),
    .B(_08907_),
    .C(_07147_),
    .Y(_07151_));
 sky130_fd_sc_hd__o311a_1 _17668_ (.A1(net301),
    .A2(_07134_),
    .A3(net300),
    .B1(_08918_),
    .C1(_07146_),
    .X(_07152_));
 sky130_fd_sc_hd__o211ai_4 _17669_ (.A1(_07134_),
    .A2(net275),
    .B1(_08918_),
    .C1(_07146_),
    .Y(_07153_));
 sky130_fd_sc_hd__a21oi_1 _17670_ (.A1(_06548_),
    .A2(_06823_),
    .B1(_06828_),
    .Y(_07155_));
 sky130_fd_sc_hd__a31o_1 _17671_ (.A1(_06548_),
    .A2(_06823_),
    .A3(_06827_),
    .B1(_06828_),
    .X(_07156_));
 sky130_fd_sc_hd__o2bb2ai_4 _17672_ (.A1_N(_07151_),
    .A2_N(_07153_),
    .B1(_07155_),
    .B2(_06825_),
    .Y(_07157_));
 sky130_fd_sc_hd__nand3_2 _17673_ (.A(_07156_),
    .B(_07153_),
    .C(_07151_),
    .Y(_07158_));
 sky130_fd_sc_hd__nand3_1 _17674_ (.A(_07157_),
    .B(_07158_),
    .C(net274),
    .Y(_07159_));
 sky130_fd_sc_hd__a31oi_4 _17675_ (.A1(_07157_),
    .A2(_07158_),
    .A3(net274),
    .B1(_07149_),
    .Y(_07160_));
 sky130_fd_sc_hd__a311oi_4 _17676_ (.A1(_07157_),
    .A2(_07158_),
    .A3(net274),
    .B1(_07149_),
    .C1(_07899_),
    .Y(_07161_));
 sky130_fd_sc_hd__a2bb2oi_2 _17677_ (.A1_N(net390),
    .A2_N(net370),
    .B1(_07150_),
    .B2(_07159_),
    .Y(_07162_));
 sky130_fd_sc_hd__inv_2 _17678_ (.A(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__o21ai_1 _17679_ (.A1(_07888_),
    .A2(_07160_),
    .B1(_06910_),
    .Y(_07164_));
 sky130_fd_sc_hd__o22ai_2 _17680_ (.A1(_06838_),
    .A2(_06909_),
    .B1(_07161_),
    .B2(_07162_),
    .Y(_07166_));
 sky130_fd_sc_hd__or3_2 _17681_ (.A(_05481_),
    .B(net269),
    .C(_07160_),
    .X(_07167_));
 sky130_fd_sc_hd__o221ai_4 _17682_ (.A1(_05481_),
    .A2(net269),
    .B1(_07161_),
    .B2(_07164_),
    .C1(_07166_),
    .Y(_07168_));
 sky130_fd_sc_hd__o21ai_1 _17683_ (.A1(_05485_),
    .A2(_07160_),
    .B1(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__a21o_1 _17684_ (.A1(_07167_),
    .A2(_07168_),
    .B1(net241),
    .X(_07170_));
 sky130_fd_sc_hd__inv_2 _17685_ (.A(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__o21ai_2 _17686_ (.A1(_06332_),
    .A2(_06845_),
    .B1(_06855_),
    .Y(_07172_));
 sky130_fd_sc_hd__o221a_1 _17687_ (.A1(_06989_),
    .A2(_07011_),
    .B1(_05485_),
    .B2(_07160_),
    .C1(_07168_),
    .X(_07173_));
 sky130_fd_sc_hd__o221ai_4 _17688_ (.A1(_06989_),
    .A2(_07011_),
    .B1(_05485_),
    .B2(_07160_),
    .C1(_07168_),
    .Y(_07174_));
 sky130_fd_sc_hd__a21oi_2 _17689_ (.A1(_07167_),
    .A2(_07168_),
    .B1(_07033_),
    .Y(_07175_));
 sky130_fd_sc_hd__o21ai_1 _17690_ (.A1(_06945_),
    .A2(_06967_),
    .B1(_07169_),
    .Y(_07177_));
 sky130_fd_sc_hd__nand3_2 _17691_ (.A(_07172_),
    .B(_07174_),
    .C(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__o21bai_2 _17692_ (.A1(_07173_),
    .A2(_07175_),
    .B1_N(_07172_),
    .Y(_07179_));
 sky130_fd_sc_hd__o211ai_2 _17693_ (.A1(net266),
    .A2(_05751_),
    .B1(_07178_),
    .C1(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__a31oi_2 _17694_ (.A1(_07179_),
    .A2(net241),
    .A3(_07178_),
    .B1(_07171_),
    .Y(_07181_));
 sky130_fd_sc_hd__a21oi_1 _17695_ (.A1(_07170_),
    .A2(_07180_),
    .B1(_05996_),
    .Y(_07182_));
 sky130_fd_sc_hd__a2bb2oi_1 _17696_ (.A1_N(_06245_),
    .A2_N(_06267_),
    .B1(_07170_),
    .B2(_07180_),
    .Y(_07183_));
 sky130_fd_sc_hd__a22o_1 _17697_ (.A1(_06256_),
    .A2(_06278_),
    .B1(_07170_),
    .B2(_07180_),
    .X(_07184_));
 sky130_fd_sc_hd__a31o_1 _17698_ (.A1(_07179_),
    .A2(net241),
    .A3(_07178_),
    .B1(_06343_),
    .X(_07185_));
 sky130_fd_sc_hd__o211a_1 _17699_ (.A1(net381),
    .A2(_06310_),
    .B1(_07170_),
    .C1(_07180_),
    .X(_07186_));
 sky130_fd_sc_hd__o21a_1 _17700_ (.A1(_06860_),
    .A2(_06864_),
    .B1(_06863_),
    .X(_07188_));
 sky130_fd_sc_hd__o21ai_2 _17701_ (.A1(_06860_),
    .A2(_06864_),
    .B1(_06863_),
    .Y(_07189_));
 sky130_fd_sc_hd__o21ai_1 _17702_ (.A1(_07183_),
    .A2(_07186_),
    .B1(_07189_),
    .Y(_07190_));
 sky130_fd_sc_hd__o211ai_2 _17703_ (.A1(_07171_),
    .A2(_07185_),
    .B1(_07188_),
    .C1(_07184_),
    .Y(_07191_));
 sky130_fd_sc_hd__a22oi_2 _17704_ (.A1(_05991_),
    .A2(_05993_),
    .B1(_07190_),
    .B2(_07191_),
    .Y(_07192_));
 sky130_fd_sc_hd__and3_1 _17705_ (.A(_07180_),
    .B(_05995_),
    .C(_07170_),
    .X(_07193_));
 sky130_fd_sc_hd__a31oi_1 _17706_ (.A1(_05996_),
    .A2(_07190_),
    .A3(_07191_),
    .B1(_07182_),
    .Y(_07194_));
 sky130_fd_sc_hd__a31o_1 _17707_ (.A1(_05996_),
    .A2(_07190_),
    .A3(_07191_),
    .B1(_07182_),
    .X(_07195_));
 sky130_fd_sc_hd__nand4_2 _17708_ (.A(_06592_),
    .B(_06595_),
    .C(_06868_),
    .D(_06869_),
    .Y(_07196_));
 sky130_fd_sc_hd__o211ai_1 _17709_ (.A1(net387),
    .A2(_06874_),
    .B1(_06883_),
    .C1(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__o2111ai_4 _17710_ (.A1(net387),
    .A2(_06874_),
    .B1(_06883_),
    .C1(_05851_),
    .D1(_07196_),
    .Y(_07199_));
 sky130_fd_sc_hd__o21ai_2 _17711_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_07197_),
    .Y(_07200_));
 sky130_fd_sc_hd__o211ai_2 _17712_ (.A1(_06291_),
    .A2(_06292_),
    .B1(_07199_),
    .C1(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__o21a_1 _17713_ (.A1(_07192_),
    .A2(_07193_),
    .B1(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__o21ai_1 _17714_ (.A1(_07192_),
    .A2(_07193_),
    .B1(_07201_),
    .Y(_07203_));
 sky130_fd_sc_hd__and4_1 _17715_ (.A(_07195_),
    .B(_07199_),
    .C(_07200_),
    .D(net212),
    .X(_07204_));
 sky130_fd_sc_hd__nand4_1 _17716_ (.A(_07195_),
    .B(_07199_),
    .C(_07200_),
    .D(net212),
    .Y(_07205_));
 sky130_fd_sc_hd__o31a_1 _17717_ (.A1(_07192_),
    .A2(_07193_),
    .A3(_07201_),
    .B1(_07203_),
    .X(_07206_));
 sky130_fd_sc_hd__nand3_2 _17718_ (.A(_06891_),
    .B(net387),
    .C(_06887_),
    .Y(_07207_));
 sky130_fd_sc_hd__o221a_2 _17719_ (.A1(_03399_),
    .A2(_05491_),
    .B1(_06886_),
    .B2(_06890_),
    .C1(net396),
    .X(_07208_));
 sky130_fd_sc_hd__o211ai_4 _17720_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_06885_),
    .C1(_06888_),
    .Y(_07210_));
 sky130_fd_sc_hd__nand3_1 _17721_ (.A(_07207_),
    .B(_07210_),
    .C(_06612_),
    .Y(_07211_));
 sky130_fd_sc_hd__o2111ai_4 _17722_ (.A1(_06608_),
    .A2(net237),
    .B1(_07207_),
    .C1(_07210_),
    .D1(_07206_),
    .Y(_07212_));
 sky130_fd_sc_hd__o21ai_2 _17723_ (.A1(_07202_),
    .A2(_07204_),
    .B1(_07211_),
    .Y(_07213_));
 sky130_fd_sc_hd__o31a_2 _17724_ (.A1(_07202_),
    .A2(_07204_),
    .A3(_07211_),
    .B1(_07213_),
    .X(_07214_));
 sky130_fd_sc_hd__o311a_1 _17725_ (.A1(_07202_),
    .A2(_07204_),
    .A3(_07211_),
    .B1(_05239_),
    .C1(_07213_),
    .X(_07215_));
 sky130_fd_sc_hd__nand3_1 _17726_ (.A(_07213_),
    .B(_05239_),
    .C(_07212_),
    .Y(_07216_));
 sky130_fd_sc_hd__a21oi_2 _17727_ (.A1(_07212_),
    .A2(_07213_),
    .B1(_05239_),
    .Y(_07217_));
 sky130_fd_sc_hd__a21o_1 _17728_ (.A1(_07212_),
    .A2(_07213_),
    .B1(_05239_),
    .X(_07218_));
 sky130_fd_sc_hd__o21ai_1 _17729_ (.A1(_07215_),
    .A2(_07217_),
    .B1(_06906_),
    .Y(_07219_));
 sky130_fd_sc_hd__a31oi_1 _17730_ (.A1(_07212_),
    .A2(_07213_),
    .A3(_05239_),
    .B1(_06906_),
    .Y(_07221_));
 sky130_fd_sc_hd__o21ai_4 _17731_ (.A1(_03289_),
    .A2(_06895_),
    .B1(_07216_),
    .Y(_07222_));
 sky130_fd_sc_hd__o211ai_4 _17732_ (.A1(_07217_),
    .A2(_07222_),
    .B1(net208),
    .C1(_07219_),
    .Y(_07223_));
 sky130_fd_sc_hd__or3_1 _17733_ (.A(net230),
    .B(_06901_),
    .C(_07214_),
    .X(_07224_));
 sky130_fd_sc_hd__o21ai_1 _17734_ (.A1(net208),
    .A2(_07214_),
    .B1(_07223_),
    .Y(_07225_));
 sky130_fd_sc_hd__or4_4 _17735_ (.A(net41),
    .B(net42),
    .C(net43),
    .D(_06285_),
    .X(_07226_));
 sky130_fd_sc_hd__and3b_4 _17736_ (.A_N(net45),
    .B(_07226_),
    .C(net409),
    .X(_07227_));
 sky130_fd_sc_hd__nand3b_4 _17737_ (.A_N(net45),
    .B(_07226_),
    .C(net409),
    .Y(_07228_));
 sky130_fd_sc_hd__a21boi_4 _17738_ (.A1(_07226_),
    .A2(net409),
    .B1_N(net45),
    .Y(_07229_));
 sky130_fd_sc_hd__a21bo_4 _17739_ (.A1(_07226_),
    .A2(net409),
    .B1_N(net45),
    .X(_07230_));
 sky130_fd_sc_hd__nor2_8 _17740_ (.A(_07227_),
    .B(net203),
    .Y(_07232_));
 sky130_fd_sc_hd__nand2_8 _17741_ (.A(_07228_),
    .B(_07230_),
    .Y(_07233_));
 sky130_fd_sc_hd__o221a_1 _17742_ (.A1(net208),
    .A2(_07214_),
    .B1(_07232_),
    .B2(_03289_),
    .C1(_07223_),
    .X(_07234_));
 sky130_fd_sc_hd__o211ai_4 _17743_ (.A1(net208),
    .A2(_07214_),
    .B1(net1),
    .C1(_07223_),
    .Y(_07235_));
 sky130_fd_sc_hd__a31oi_2 _17744_ (.A1(net1),
    .A2(_07225_),
    .A3(net185),
    .B1(_07234_),
    .Y(_07236_));
 sky130_fd_sc_hd__or3_1 _17745_ (.A(_05051_),
    .B(_06908_),
    .C(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__o21ai_1 _17746_ (.A1(_05051_),
    .A2(_06908_),
    .B1(_07236_),
    .Y(_07238_));
 sky130_fd_sc_hd__and2_1 _17747_ (.A(_07237_),
    .B(_07238_),
    .X(net77));
 sky130_fd_sc_hd__o2bb2a_1 _17748_ (.A1_N(_06908_),
    .A2_N(_07236_),
    .B1(_04832_),
    .B2(_04942_),
    .X(_07239_));
 sky130_fd_sc_hd__or4_4 _17749_ (.A(net10),
    .B(net11),
    .C(net13),
    .D(_06304_),
    .X(_07240_));
 sky130_fd_sc_hd__and3b_4 _17750_ (.A_N(net14),
    .B(_07240_),
    .C(net410),
    .X(_07242_));
 sky130_fd_sc_hd__a21boi_4 _17751_ (.A1(_07240_),
    .A2(net410),
    .B1_N(net14),
    .Y(_07243_));
 sky130_fd_sc_hd__and3_4 _17752_ (.A(_07240_),
    .B(net14),
    .C(net410),
    .X(_07244_));
 sky130_fd_sc_hd__a21oi_4 _17753_ (.A1(_07240_),
    .A2(net410),
    .B1(net14),
    .Y(_07245_));
 sky130_fd_sc_hd__nor2_8 _17754_ (.A(_07242_),
    .B(net248),
    .Y(_07246_));
 sky130_fd_sc_hd__nor2_8 _17755_ (.A(_07244_),
    .B(net247),
    .Y(_07247_));
 sky130_fd_sc_hd__o21a_1 _17756_ (.A1(_07242_),
    .A2(_07243_),
    .B1(net33),
    .X(_07248_));
 sky130_fd_sc_hd__or3_4 _17757_ (.A(_07245_),
    .B(_03178_),
    .C(_07244_),
    .X(_07249_));
 sky130_fd_sc_hd__or4_1 _17758_ (.A(_03178_),
    .B(_06918_),
    .C(_06920_),
    .D(net224),
    .X(_07250_));
 sky130_fd_sc_hd__or3_1 _17759_ (.A(_06914_),
    .B(_06916_),
    .C(_07248_),
    .X(_07251_));
 sky130_fd_sc_hd__o21ai_4 _17760_ (.A1(_06925_),
    .A2(net224),
    .B1(_07251_),
    .Y(_07253_));
 sky130_fd_sc_hd__a31oi_4 _17761_ (.A1(_06633_),
    .A2(_06931_),
    .A3(_06930_),
    .B1(_06927_),
    .Y(_07254_));
 sky130_fd_sc_hd__a31o_2 _17762_ (.A1(_06633_),
    .A2(_06931_),
    .A3(_06930_),
    .B1(_06927_),
    .X(_07255_));
 sky130_fd_sc_hd__a21oi_2 _17763_ (.A1(_06928_),
    .A2(_06933_),
    .B1(_07253_),
    .Y(_07256_));
 sky130_fd_sc_hd__a21o_1 _17764_ (.A1(_06928_),
    .A2(_06933_),
    .B1(_07253_),
    .X(_07257_));
 sky130_fd_sc_hd__nand2_1 _17765_ (.A(_07254_),
    .B(_07253_),
    .Y(_07258_));
 sky130_fd_sc_hd__a21oi_4 _17766_ (.A1(_07257_),
    .A2(_07258_),
    .B1(_05185_),
    .Y(_07259_));
 sky130_fd_sc_hd__a31o_1 _17767_ (.A1(_06928_),
    .A2(_06933_),
    .A3(_07253_),
    .B1(_05185_),
    .X(_07260_));
 sky130_fd_sc_hd__a211o_2 _17768_ (.A1(_05185_),
    .A2(_07249_),
    .B1(net388),
    .C1(_07259_),
    .X(_07261_));
 sky130_fd_sc_hd__o221a_1 _17769_ (.A1(net405),
    .A2(_07249_),
    .B1(_07256_),
    .B2(_07260_),
    .C1(net234),
    .X(_07262_));
 sky130_fd_sc_hd__o221ai_4 _17770_ (.A1(net405),
    .A2(_07249_),
    .B1(_07256_),
    .B2(_07260_),
    .C1(net234),
    .Y(_07264_));
 sky130_fd_sc_hd__a22o_2 _17771_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_07249_),
    .B2(_05185_),
    .X(_07265_));
 sky130_fd_sc_hd__o21a_2 _17772_ (.A1(_07265_),
    .A2(_07259_),
    .B1(_07264_),
    .X(_07266_));
 sky130_fd_sc_hd__o21ai_2 _17773_ (.A1(_07265_),
    .A2(_07259_),
    .B1(_07264_),
    .Y(_07267_));
 sky130_fd_sc_hd__o22ai_4 _17774_ (.A1(_06935_),
    .A2(_06943_),
    .B1(_06947_),
    .B2(_06940_),
    .Y(_07268_));
 sky130_fd_sc_hd__nand2_1 _17775_ (.A(_07268_),
    .B(_07266_),
    .Y(_07269_));
 sky130_fd_sc_hd__o21ai_1 _17776_ (.A1(_06314_),
    .A2(_06939_),
    .B1(_07267_),
    .Y(_07270_));
 sky130_fd_sc_hd__o211ai_2 _17777_ (.A1(_06947_),
    .A2(_06940_),
    .B1(_06946_),
    .C1(_07267_),
    .Y(_07271_));
 sky130_fd_sc_hd__a21oi_2 _17778_ (.A1(_07268_),
    .A2(_07266_),
    .B1(_05392_),
    .Y(_07272_));
 sky130_fd_sc_hd__o211ai_4 _17779_ (.A1(_07270_),
    .A2(_06949_),
    .B1(net388),
    .C1(_07269_),
    .Y(_07273_));
 sky130_fd_sc_hd__a21boi_4 _17780_ (.A1(_07272_),
    .A2(_07271_),
    .B1_N(_07261_),
    .Y(_07275_));
 sky130_fd_sc_hd__nand2_1 _17781_ (.A(_07261_),
    .B(_07273_),
    .Y(_07276_));
 sky130_fd_sc_hd__a2bb2oi_4 _17782_ (.A1_N(_06305_),
    .A2_N(net283),
    .B1(_07261_),
    .B2(_07273_),
    .Y(_07277_));
 sky130_fd_sc_hd__a21oi_1 _17783_ (.A1(_07272_),
    .A2(_07271_),
    .B1(net251),
    .Y(_07278_));
 sky130_fd_sc_hd__and3_2 _17784_ (.A(_07273_),
    .B(_06314_),
    .C(_07261_),
    .X(_07279_));
 sky130_fd_sc_hd__a21oi_1 _17785_ (.A1(_07261_),
    .A2(_07278_),
    .B1(_07277_),
    .Y(_07280_));
 sky130_fd_sc_hd__o32ai_1 _17786_ (.A1(net286),
    .A2(_06012_),
    .A3(_06953_),
    .B1(_06959_),
    .B2(_06960_),
    .Y(_07281_));
 sky130_fd_sc_hd__o22ai_1 _17787_ (.A1(_06959_),
    .A2(_06960_),
    .B1(_07277_),
    .B2(_07279_),
    .Y(_07282_));
 sky130_fd_sc_hd__o221ai_4 _17788_ (.A1(_06959_),
    .A2(_06960_),
    .B1(_07277_),
    .B2(_07279_),
    .C1(_06955_),
    .Y(_07283_));
 sky130_fd_sc_hd__nand2_1 _17789_ (.A(_07281_),
    .B(_07280_),
    .Y(_07284_));
 sky130_fd_sc_hd__and3_1 _17790_ (.A(_05687_),
    .B(_05709_),
    .C(_07276_),
    .X(_07286_));
 sky130_fd_sc_hd__or3_1 _17791_ (.A(net384),
    .B(net383),
    .C(_07275_),
    .X(_07287_));
 sky130_fd_sc_hd__o221a_1 _17792_ (.A1(net384),
    .A2(net383),
    .B1(_06957_),
    .B2(_07282_),
    .C1(_07284_),
    .X(_07288_));
 sky130_fd_sc_hd__nand3_2 _17793_ (.A(_07284_),
    .B(net359),
    .C(_07283_),
    .Y(_07289_));
 sky130_fd_sc_hd__o31a_4 _17794_ (.A1(net384),
    .A2(net383),
    .A3(_07275_),
    .B1(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__or3_1 _17795_ (.A(_06793_),
    .B(_06815_),
    .C(_07290_),
    .X(_07291_));
 sky130_fd_sc_hd__a2bb2oi_2 _17796_ (.A1_N(_06009_),
    .A2_N(_06010_),
    .B1(_07287_),
    .B2(_07289_),
    .Y(_07292_));
 sky130_fd_sc_hd__o22ai_2 _17797_ (.A1(_06009_),
    .A2(_06010_),
    .B1(_07286_),
    .B2(_07288_),
    .Y(_07293_));
 sky130_fd_sc_hd__a31oi_1 _17798_ (.A1(_07284_),
    .A2(net359),
    .A3(_07283_),
    .B1(net253),
    .Y(_07294_));
 sky130_fd_sc_hd__a31o_1 _17799_ (.A1(_07284_),
    .A2(net359),
    .A3(_07283_),
    .B1(net253),
    .X(_07295_));
 sky130_fd_sc_hd__o221a_1 _17800_ (.A1(net286),
    .A2(_06012_),
    .B1(_07275_),
    .B2(net359),
    .C1(_07289_),
    .X(_07297_));
 sky130_fd_sc_hd__a21oi_2 _17801_ (.A1(_07287_),
    .A2(_07294_),
    .B1(_07292_),
    .Y(_07298_));
 sky130_fd_sc_hd__o21ai_2 _17802_ (.A1(_07286_),
    .A2(_07295_),
    .B1(_07293_),
    .Y(_07299_));
 sky130_fd_sc_hd__o31a_1 _17803_ (.A1(_06977_),
    .A2(_06686_),
    .A3(_06684_),
    .B1(_06971_),
    .X(_07300_));
 sky130_fd_sc_hd__a21oi_2 _17804_ (.A1(_07300_),
    .A2(_06985_),
    .B1(_06966_),
    .Y(_07301_));
 sky130_fd_sc_hd__o221ai_4 _17805_ (.A1(_06969_),
    .A2(_06954_),
    .B1(_06966_),
    .B2(_06986_),
    .C1(_07298_),
    .Y(_07302_));
 sky130_fd_sc_hd__o221ai_4 _17806_ (.A1(_07292_),
    .A2(_07297_),
    .B1(_06973_),
    .B2(_06987_),
    .C1(_06968_),
    .Y(_07303_));
 sky130_fd_sc_hd__nand3_4 _17807_ (.A(_07302_),
    .B(_07303_),
    .C(net357),
    .Y(_07304_));
 sky130_fd_sc_hd__o21ai_2 _17808_ (.A1(net357),
    .A2(_07290_),
    .B1(_07304_),
    .Y(_07305_));
 sky130_fd_sc_hd__a2bb2oi_2 _17809_ (.A1_N(_05760_),
    .A2_N(net290),
    .B1(_07291_),
    .B2(_07304_),
    .Y(_07306_));
 sky130_fd_sc_hd__a22o_1 _17810_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_07291_),
    .B2(_07304_),
    .X(_07308_));
 sky130_fd_sc_hd__o221a_1 _17811_ (.A1(_05765_),
    .A2(net289),
    .B1(_07290_),
    .B2(net357),
    .C1(_07304_),
    .X(_07309_));
 sky130_fd_sc_hd__o221ai_4 _17812_ (.A1(_05765_),
    .A2(net289),
    .B1(_07290_),
    .B2(net357),
    .C1(_07304_),
    .Y(_07310_));
 sky130_fd_sc_hd__nor2_1 _17813_ (.A(_07306_),
    .B(_07309_),
    .Y(_07311_));
 sky130_fd_sc_hd__a22oi_2 _17814_ (.A1(_06965_),
    .A2(_07003_),
    .B1(_07007_),
    .B2(_07010_),
    .Y(_07312_));
 sky130_fd_sc_hd__o22ai_4 _17815_ (.A1(_07004_),
    .A2(_06964_),
    .B1(_07009_),
    .B2(_07006_),
    .Y(_07313_));
 sky130_fd_sc_hd__nand3_1 _17816_ (.A(_07308_),
    .B(_07310_),
    .C(_07313_),
    .Y(_07314_));
 sky130_fd_sc_hd__o21ai_1 _17817_ (.A1(_07306_),
    .A2(_07309_),
    .B1(_07312_),
    .Y(_07315_));
 sky130_fd_sc_hd__nand3_1 _17818_ (.A(_07308_),
    .B(_07310_),
    .C(_07312_),
    .Y(_07316_));
 sky130_fd_sc_hd__o21ai_1 _17819_ (.A1(_07306_),
    .A2(_07309_),
    .B1(_07313_),
    .Y(_07317_));
 sky130_fd_sc_hd__nand3_2 _17820_ (.A(_07315_),
    .B(net355),
    .C(_07314_),
    .Y(_07319_));
 sky130_fd_sc_hd__a211o_1 _17821_ (.A1(_07291_),
    .A2(_07304_),
    .B1(net373),
    .C1(net371),
    .X(_07320_));
 sky130_fd_sc_hd__o211ai_4 _17822_ (.A1(net373),
    .A2(net371),
    .B1(_07316_),
    .C1(_07317_),
    .Y(_07321_));
 sky130_fd_sc_hd__o21a_1 _17823_ (.A1(net355),
    .A2(_07305_),
    .B1(_07319_),
    .X(_07322_));
 sky130_fd_sc_hd__and3_1 _17824_ (.A(_07322_),
    .B(_08711_),
    .C(_08689_),
    .X(_07323_));
 sky130_fd_sc_hd__a211o_1 _17825_ (.A1(_07320_),
    .A2(_07321_),
    .B1(net353),
    .C1(net352),
    .X(_07324_));
 sky130_fd_sc_hd__o211a_1 _17826_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_07320_),
    .C1(_07321_),
    .X(_07325_));
 sky130_fd_sc_hd__o211ai_4 _17827_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_07320_),
    .C1(_07321_),
    .Y(_07326_));
 sky130_fd_sc_hd__o211ai_4 _17828_ (.A1(_07305_),
    .A2(net355),
    .B1(net291),
    .C1(_07319_),
    .Y(_07327_));
 sky130_fd_sc_hd__nand2_1 _17829_ (.A(_07326_),
    .B(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__nand2_1 _17830_ (.A(_07027_),
    .B(_07020_),
    .Y(_07330_));
 sky130_fd_sc_hd__o22ai_4 _17831_ (.A1(_07001_),
    .A2(_07023_),
    .B1(_07019_),
    .B2(_07028_),
    .Y(_07331_));
 sky130_fd_sc_hd__a22oi_1 _17832_ (.A1(_07326_),
    .A2(_07327_),
    .B1(_07330_),
    .B2(_07025_),
    .Y(_07332_));
 sky130_fd_sc_hd__nand2_2 _17833_ (.A(_07328_),
    .B(_07331_),
    .Y(_07333_));
 sky130_fd_sc_hd__o2111a_1 _17834_ (.A1(net293),
    .A2(_07018_),
    .B1(_07326_),
    .C1(_07327_),
    .D1(_07330_),
    .X(_07334_));
 sky130_fd_sc_hd__o2111ai_4 _17835_ (.A1(net293),
    .A2(_07018_),
    .B1(_07326_),
    .C1(_07327_),
    .D1(_07330_),
    .Y(_07335_));
 sky130_fd_sc_hd__nand3_2 _17836_ (.A(_07333_),
    .B(_07335_),
    .C(net338),
    .Y(_07336_));
 sky130_fd_sc_hd__o22ai_2 _17837_ (.A1(net353),
    .A2(net352),
    .B1(_07332_),
    .B2(_07334_),
    .Y(_07337_));
 sky130_fd_sc_hd__a31o_1 _17838_ (.A1(_07333_),
    .A2(_07335_),
    .A3(net338),
    .B1(_07323_),
    .X(_07338_));
 sky130_fd_sc_hd__o21a_1 _17839_ (.A1(net299),
    .A2(_07039_),
    .B1(_07046_),
    .X(_07339_));
 sky130_fd_sc_hd__o21ai_1 _17840_ (.A1(_07046_),
    .A2(_07042_),
    .B1(_07041_),
    .Y(_07341_));
 sky130_fd_sc_hd__a21oi_1 _17841_ (.A1(_07045_),
    .A2(_07043_),
    .B1(_07040_),
    .Y(_07342_));
 sky130_fd_sc_hd__a311oi_4 _17842_ (.A1(_07333_),
    .A2(_07335_),
    .A3(net338),
    .B1(net293),
    .C1(_07323_),
    .Y(_07343_));
 sky130_fd_sc_hd__nand4_2 _17843_ (.A(_05243_),
    .B(_05245_),
    .C(_07324_),
    .D(_07336_),
    .Y(_07344_));
 sky130_fd_sc_hd__a2bb2oi_2 _17844_ (.A1_N(_05242_),
    .A2_N(net314),
    .B1(_07324_),
    .B2(_07336_),
    .Y(_07345_));
 sky130_fd_sc_hd__o221ai_4 _17845_ (.A1(_05242_),
    .A2(net314),
    .B1(_07322_),
    .B2(net338),
    .C1(_07337_),
    .Y(_07346_));
 sky130_fd_sc_hd__nand3_1 _17846_ (.A(_07342_),
    .B(_07344_),
    .C(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__o2bb2ai_1 _17847_ (.A1_N(_07041_),
    .A2_N(_07053_),
    .B1(_07343_),
    .B2(_07345_),
    .Y(_07348_));
 sky130_fd_sc_hd__nand3_1 _17848_ (.A(_07348_),
    .B(net336),
    .C(_07347_),
    .Y(_07349_));
 sky130_fd_sc_hd__a211o_1 _17849_ (.A1(_07324_),
    .A2(_07336_),
    .B1(_09785_),
    .C1(net349),
    .X(_07350_));
 sky130_fd_sc_hd__inv_2 _17850_ (.A(_07350_),
    .Y(_07352_));
 sky130_fd_sc_hd__nand3_1 _17851_ (.A(_07346_),
    .B(_07341_),
    .C(_07344_),
    .Y(_07353_));
 sky130_fd_sc_hd__o22ai_2 _17852_ (.A1(_07042_),
    .A2(_07339_),
    .B1(_07343_),
    .B2(_07345_),
    .Y(_07354_));
 sky130_fd_sc_hd__o211ai_2 _17853_ (.A1(_09785_),
    .A2(net349),
    .B1(_07353_),
    .C1(_07354_),
    .Y(_07355_));
 sky130_fd_sc_hd__a31o_1 _17854_ (.A1(net336),
    .A2(_07353_),
    .A3(_07354_),
    .B1(_07352_),
    .X(_07356_));
 sky130_fd_sc_hd__inv_2 _17855_ (.A(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__o211a_1 _17856_ (.A1(_07338_),
    .A2(net336),
    .B1(net298),
    .C1(_07349_),
    .X(_07358_));
 sky130_fd_sc_hd__o211ai_4 _17857_ (.A1(_07338_),
    .A2(net336),
    .B1(net298),
    .C1(_07349_),
    .Y(_07359_));
 sky130_fd_sc_hd__a31o_1 _17858_ (.A1(_07354_),
    .A2(net336),
    .A3(_07353_),
    .B1(net298),
    .X(_07360_));
 sky130_fd_sc_hd__and3_1 _17859_ (.A(_07355_),
    .B(net299),
    .C(_07350_),
    .X(_07361_));
 sky130_fd_sc_hd__nand3_1 _17860_ (.A(_07355_),
    .B(net299),
    .C(_07350_),
    .Y(_07363_));
 sky130_fd_sc_hd__nand2_2 _17861_ (.A(_07359_),
    .B(_07363_),
    .Y(_07364_));
 sky130_fd_sc_hd__a31oi_4 _17862_ (.A1(_07062_),
    .A2(_07069_),
    .A3(_07071_),
    .B1(_07058_),
    .Y(_07365_));
 sky130_fd_sc_hd__o22ai_1 _17863_ (.A1(_02137_),
    .A2(_07056_),
    .B1(_07068_),
    .B2(_07079_),
    .Y(_07366_));
 sky130_fd_sc_hd__a21oi_4 _17864_ (.A1(_07059_),
    .A2(_07080_),
    .B1(_07364_),
    .Y(_07367_));
 sky130_fd_sc_hd__o211ai_1 _17865_ (.A1(_07360_),
    .A2(_07352_),
    .B1(_07359_),
    .C1(_07366_),
    .Y(_07368_));
 sky130_fd_sc_hd__nand2_1 _17866_ (.A(_07365_),
    .B(_07364_),
    .Y(_07369_));
 sky130_fd_sc_hd__o2bb2ai_4 _17867_ (.A1_N(_07364_),
    .A2_N(_07365_),
    .B1(net347),
    .B2(net346),
    .Y(_07370_));
 sky130_fd_sc_hd__nand3_2 _17868_ (.A(_07368_),
    .B(_07369_),
    .C(net334),
    .Y(_07371_));
 sky130_fd_sc_hd__a211o_1 _17869_ (.A1(_07350_),
    .A2(_07355_),
    .B1(net347),
    .C1(net346),
    .X(_07372_));
 sky130_fd_sc_hd__o22ai_4 _17870_ (.A1(net334),
    .A2(_07357_),
    .B1(_07367_),
    .B2(_07370_),
    .Y(_07374_));
 sky130_fd_sc_hd__o22a_1 _17871_ (.A1(_06757_),
    .A2(_07092_),
    .B1(net320),
    .B2(_07084_),
    .X(_07375_));
 sky130_fd_sc_hd__o21ai_1 _17872_ (.A1(_06757_),
    .A2(_07092_),
    .B1(_07091_),
    .Y(_07376_));
 sky130_fd_sc_hd__a22oi_4 _17873_ (.A1(_07078_),
    .A2(_07087_),
    .B1(_07091_),
    .B2(_07094_),
    .Y(_07377_));
 sky130_fd_sc_hd__a31o_1 _17874_ (.A1(net320),
    .A2(_07078_),
    .A3(_07083_),
    .B1(_07375_),
    .X(_07378_));
 sky130_fd_sc_hd__a22oi_4 _17875_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_07371_),
    .B2(_07372_),
    .Y(_07379_));
 sky130_fd_sc_hd__o21ai_2 _17876_ (.A1(_02049_),
    .A2(net342),
    .B1(_07374_),
    .Y(_07380_));
 sky130_fd_sc_hd__o221a_2 _17877_ (.A1(net334),
    .A2(_07357_),
    .B1(_07367_),
    .B2(_07370_),
    .C1(_02137_),
    .X(_07381_));
 sky130_fd_sc_hd__o221ai_4 _17878_ (.A1(net334),
    .A2(_07357_),
    .B1(_07367_),
    .B2(_07370_),
    .C1(_02137_),
    .Y(_07382_));
 sky130_fd_sc_hd__o211ai_1 _17879_ (.A1(_07089_),
    .A2(_07375_),
    .B1(_07380_),
    .C1(_07382_),
    .Y(_07383_));
 sky130_fd_sc_hd__o21ai_1 _17880_ (.A1(_07379_),
    .A2(_07381_),
    .B1(_07377_),
    .Y(_07385_));
 sky130_fd_sc_hd__o22ai_4 _17881_ (.A1(_07089_),
    .A2(_07375_),
    .B1(_07379_),
    .B2(_07381_),
    .Y(_07386_));
 sky130_fd_sc_hd__nand3_2 _17882_ (.A(_07380_),
    .B(_07382_),
    .C(_07377_),
    .Y(_07387_));
 sky130_fd_sc_hd__nand3_2 _17883_ (.A(_07385_),
    .B(net312),
    .C(_07383_),
    .Y(_07388_));
 sky130_fd_sc_hd__a21oi_1 _17884_ (.A1(_07371_),
    .A2(_07372_),
    .B1(net312),
    .Y(_07389_));
 sky130_fd_sc_hd__a211o_1 _17885_ (.A1(_07371_),
    .A2(_07372_),
    .B1(_12670_),
    .C1(_12681_),
    .X(_07390_));
 sky130_fd_sc_hd__nand3_2 _17886_ (.A(_07386_),
    .B(_07387_),
    .C(net312),
    .Y(_07391_));
 sky130_fd_sc_hd__o211a_2 _17887_ (.A1(_07374_),
    .A2(net312),
    .B1(_00066_),
    .C1(_07388_),
    .X(_07392_));
 sky130_fd_sc_hd__a211o_1 _17888_ (.A1(_07390_),
    .A2(_07391_),
    .B1(net324),
    .C1(_00033_),
    .X(_07393_));
 sky130_fd_sc_hd__a311oi_4 _17889_ (.A1(_07386_),
    .A2(_07387_),
    .A3(net312),
    .B1(_07389_),
    .C1(net319),
    .Y(_07394_));
 sky130_fd_sc_hd__nand3_4 _17890_ (.A(_07391_),
    .B(net320),
    .C(_07390_),
    .Y(_07396_));
 sky130_fd_sc_hd__a2bb2oi_1 _17891_ (.A1_N(_00174_),
    .A2_N(_00196_),
    .B1(_07390_),
    .B2(_07391_),
    .Y(_07397_));
 sky130_fd_sc_hd__o211ai_4 _17892_ (.A1(_07374_),
    .A2(net312),
    .B1(net319),
    .C1(_07388_),
    .Y(_07398_));
 sky130_fd_sc_hd__a21oi_1 _17893_ (.A1(net325),
    .A2(_07103_),
    .B1(_07106_),
    .Y(_07399_));
 sky130_fd_sc_hd__o21ai_1 _17894_ (.A1(_06773_),
    .A2(_07104_),
    .B1(_07111_),
    .Y(_07400_));
 sky130_fd_sc_hd__a21oi_2 _17895_ (.A1(_07108_),
    .A2(_07106_),
    .B1(_07109_),
    .Y(_07401_));
 sky130_fd_sc_hd__o2bb2ai_4 _17896_ (.A1_N(_07396_),
    .A2_N(_07398_),
    .B1(_07399_),
    .B2(_07107_),
    .Y(_07402_));
 sky130_fd_sc_hd__o2111ai_4 _17897_ (.A1(net325),
    .A2(_07103_),
    .B1(_07396_),
    .C1(_07398_),
    .D1(_07400_),
    .Y(_07403_));
 sky130_fd_sc_hd__nand3_1 _17898_ (.A(_07402_),
    .B(_07403_),
    .C(net309),
    .Y(_07404_));
 sky130_fd_sc_hd__a31oi_4 _17899_ (.A1(_07402_),
    .A2(_07403_),
    .A3(net309),
    .B1(_07392_),
    .Y(_07405_));
 sky130_fd_sc_hd__a311o_1 _17900_ (.A1(_07402_),
    .A2(_07403_),
    .A3(net309),
    .B1(_01962_),
    .C1(_07392_),
    .X(_07407_));
 sky130_fd_sc_hd__a21oi_2 _17901_ (.A1(_07120_),
    .A2(net330),
    .B1(_07127_),
    .Y(_07408_));
 sky130_fd_sc_hd__a311oi_4 _17902_ (.A1(_07402_),
    .A2(_07403_),
    .A3(net309),
    .B1(_07392_),
    .C1(net325),
    .Y(_07409_));
 sky130_fd_sc_hd__a311o_1 _17903_ (.A1(_07402_),
    .A2(_07403_),
    .A3(net309),
    .B1(_07392_),
    .C1(net325),
    .X(_07410_));
 sky130_fd_sc_hd__a2bb2oi_1 _17904_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_07393_),
    .B2(_07404_),
    .Y(_07411_));
 sky130_fd_sc_hd__a2bb2o_1 _17905_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_07393_),
    .B2(_07404_),
    .X(_07412_));
 sky130_fd_sc_hd__o211ai_1 _17906_ (.A1(_07124_),
    .A2(_07408_),
    .B1(_07410_),
    .C1(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__o2bb2ai_1 _17907_ (.A1_N(_07123_),
    .A2_N(_07129_),
    .B1(_07409_),
    .B2(_07411_),
    .Y(_07414_));
 sky130_fd_sc_hd__nand3_1 _17908_ (.A(_07413_),
    .B(_07414_),
    .C(_01962_),
    .Y(_07415_));
 sky130_fd_sc_hd__or3_1 _17909_ (.A(net306),
    .B(net303),
    .C(_07405_),
    .X(_07416_));
 sky130_fd_sc_hd__o2bb2ai_1 _17910_ (.A1_N(_07123_),
    .A2_N(_07129_),
    .B1(_07405_),
    .B2(_12888_),
    .Y(_07418_));
 sky130_fd_sc_hd__o22ai_2 _17911_ (.A1(_07124_),
    .A2(_07408_),
    .B1(_07409_),
    .B2(_07411_),
    .Y(_07419_));
 sky130_fd_sc_hd__o221ai_4 _17912_ (.A1(net306),
    .A2(net303),
    .B1(_07409_),
    .B2(_07418_),
    .C1(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__o21ai_2 _17913_ (.A1(net280),
    .A2(_07405_),
    .B1(_07420_),
    .Y(_07421_));
 sky130_fd_sc_hd__o211ai_4 _17914_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_07407_),
    .C1(_07415_),
    .Y(_07422_));
 sky130_fd_sc_hd__inv_2 _17915_ (.A(_07422_),
    .Y(_07423_));
 sky130_fd_sc_hd__and3_1 _17916_ (.A(_07420_),
    .B(net331),
    .C(_07416_),
    .X(_07424_));
 sky130_fd_sc_hd__o211ai_4 _17917_ (.A1(net280),
    .A2(_07405_),
    .B1(net331),
    .C1(_07420_),
    .Y(_07425_));
 sky130_fd_sc_hd__a21oi_1 _17918_ (.A1(net348),
    .A2(_07134_),
    .B1(_07140_),
    .Y(_07426_));
 sky130_fd_sc_hd__o32a_1 _17919_ (.A1(_09927_),
    .A2(_09949_),
    .A3(_07134_),
    .B1(_07140_),
    .B2(_07135_),
    .X(_07427_));
 sky130_fd_sc_hd__a21oi_1 _17920_ (.A1(_07138_),
    .A2(_07140_),
    .B1(_07135_),
    .Y(_07429_));
 sky130_fd_sc_hd__o2111ai_4 _17921_ (.A1(_07137_),
    .A2(_07139_),
    .B1(_07422_),
    .C1(_07425_),
    .D1(_07136_),
    .Y(_07430_));
 sky130_fd_sc_hd__a21o_1 _17922_ (.A1(_07422_),
    .A2(_07425_),
    .B1(_07429_),
    .X(_07431_));
 sky130_fd_sc_hd__o211ai_4 _17923_ (.A1(net301),
    .A2(net300),
    .B1(_07430_),
    .C1(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__a2bb2o_2 _17924_ (.A1_N(_03986_),
    .A2_N(_03997_),
    .B1(_07416_),
    .B2(_07420_),
    .X(_07433_));
 sky130_fd_sc_hd__inv_2 _17925_ (.A(_07433_),
    .Y(_07434_));
 sky130_fd_sc_hd__o2bb2ai_2 _17926_ (.A1_N(_07422_),
    .A2_N(_07425_),
    .B1(_07426_),
    .B2(_07137_),
    .Y(_07435_));
 sky130_fd_sc_hd__and3_1 _17927_ (.A(_07427_),
    .B(_07425_),
    .C(_07422_),
    .X(_07436_));
 sky130_fd_sc_hd__nand3_4 _17928_ (.A(_07427_),
    .B(_07425_),
    .C(_07422_),
    .Y(_07437_));
 sky130_fd_sc_hd__nand3_2 _17929_ (.A(_07435_),
    .B(_07437_),
    .C(net275),
    .Y(_07438_));
 sky130_fd_sc_hd__a31oi_4 _17930_ (.A1(_07435_),
    .A2(_07437_),
    .A3(net275),
    .B1(_07434_),
    .Y(_07440_));
 sky130_fd_sc_hd__a311o_1 _17931_ (.A1(_07435_),
    .A2(_07437_),
    .A3(net275),
    .B1(_05233_),
    .C1(_07434_),
    .X(_07441_));
 sky130_fd_sc_hd__a2bb2oi_2 _17932_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_07433_),
    .B2(_07438_),
    .Y(_07442_));
 sky130_fd_sc_hd__o211ai_4 _17933_ (.A1(net275),
    .A2(_07421_),
    .B1(_07432_),
    .C1(net348),
    .Y(_07443_));
 sky130_fd_sc_hd__o211a_2 _17934_ (.A1(_09971_),
    .A2(_09993_),
    .B1(_07433_),
    .C1(_07438_),
    .X(_07444_));
 sky130_fd_sc_hd__o211ai_2 _17935_ (.A1(_09971_),
    .A2(_09993_),
    .B1(_07433_),
    .C1(_07438_),
    .Y(_07445_));
 sky130_fd_sc_hd__a32oi_2 _17936_ (.A1(_07148_),
    .A2(_08907_),
    .A3(_07147_),
    .B1(_06829_),
    .B2(_06830_),
    .Y(_07446_));
 sky130_fd_sc_hd__a21oi_2 _17937_ (.A1(_07156_),
    .A2(_07151_),
    .B1(_07152_),
    .Y(_07447_));
 sky130_fd_sc_hd__o21ai_2 _17938_ (.A1(_07442_),
    .A2(_07444_),
    .B1(_07447_),
    .Y(_07448_));
 sky130_fd_sc_hd__o2bb2a_1 _17939_ (.A1_N(_10015_),
    .A2_N(_07440_),
    .B1(_07446_),
    .B2(_07152_),
    .X(_07449_));
 sky130_fd_sc_hd__o211ai_2 _17940_ (.A1(_07152_),
    .A2(_07446_),
    .B1(_07445_),
    .C1(_07443_),
    .Y(_07451_));
 sky130_fd_sc_hd__nand3_1 _17941_ (.A(_07447_),
    .B(_07445_),
    .C(_07443_),
    .Y(_07452_));
 sky130_fd_sc_hd__a21o_1 _17942_ (.A1(_07443_),
    .A2(_07445_),
    .B1(_07447_),
    .X(_07453_));
 sky130_fd_sc_hd__o211ai_1 _17943_ (.A1(net297),
    .A2(_05232_),
    .B1(_07452_),
    .C1(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__o211a_1 _17944_ (.A1(net275),
    .A2(_07421_),
    .B1(_07432_),
    .C1(_05234_),
    .X(_07455_));
 sky130_fd_sc_hd__inv_2 _17945_ (.A(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__nand3_2 _17946_ (.A(_07448_),
    .B(_07451_),
    .C(net274),
    .Y(_07457_));
 sky130_fd_sc_hd__o31a_1 _17947_ (.A1(net297),
    .A2(_05232_),
    .A3(_07440_),
    .B1(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__a311o_1 _17948_ (.A1(_07448_),
    .A2(_07451_),
    .A3(_05233_),
    .B1(_07455_),
    .C1(_05485_),
    .X(_07459_));
 sky130_fd_sc_hd__o31a_1 _17949_ (.A1(net369),
    .A2(_07866_),
    .A3(_07160_),
    .B1(_06911_),
    .X(_07460_));
 sky130_fd_sc_hd__a21oi_1 _17950_ (.A1(_07888_),
    .A2(_07160_),
    .B1(_06911_),
    .Y(_07462_));
 sky130_fd_sc_hd__o21bai_2 _17951_ (.A1(_06911_),
    .A2(_07161_),
    .B1_N(_07162_),
    .Y(_07463_));
 sky130_fd_sc_hd__a311oi_2 _17952_ (.A1(_07448_),
    .A2(_07451_),
    .A3(_05233_),
    .B1(_07455_),
    .C1(_08918_),
    .Y(_07464_));
 sky130_fd_sc_hd__o211ai_4 _17953_ (.A1(net274),
    .A2(_07440_),
    .B1(_08907_),
    .C1(_07457_),
    .Y(_07465_));
 sky130_fd_sc_hd__a2bb2oi_2 _17954_ (.A1_N(_08819_),
    .A2_N(net367),
    .B1(_07456_),
    .B2(_07457_),
    .Y(_07466_));
 sky130_fd_sc_hd__o211ai_1 _17955_ (.A1(_08819_),
    .A2(net367),
    .B1(_07441_),
    .C1(_07454_),
    .Y(_07467_));
 sky130_fd_sc_hd__o2111ai_1 _17956_ (.A1(_06911_),
    .A2(_07161_),
    .B1(_07163_),
    .C1(_07465_),
    .D1(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__o22ai_1 _17957_ (.A1(_07162_),
    .A2(_07462_),
    .B1(_07464_),
    .B2(_07466_),
    .Y(_07469_));
 sky130_fd_sc_hd__nand3_1 _17958_ (.A(_07469_),
    .B(_05485_),
    .C(_07468_),
    .Y(_07470_));
 sky130_fd_sc_hd__o211ai_1 _17959_ (.A1(_07162_),
    .A2(_07462_),
    .B1(_07465_),
    .C1(_07467_),
    .Y(_07471_));
 sky130_fd_sc_hd__o22ai_1 _17960_ (.A1(_07161_),
    .A2(_07460_),
    .B1(_07464_),
    .B2(_07466_),
    .Y(_07473_));
 sky130_fd_sc_hd__nand3_2 _17961_ (.A(_07473_),
    .B(_05485_),
    .C(_07471_),
    .Y(_07474_));
 sky130_fd_sc_hd__o31a_2 _17962_ (.A1(_05481_),
    .A2(net269),
    .A3(_07458_),
    .B1(_07474_),
    .X(_07475_));
 sky130_fd_sc_hd__and3_1 _17963_ (.A(_05754_),
    .B(_07459_),
    .C(_07470_),
    .X(_07476_));
 sky130_fd_sc_hd__or2_1 _17964_ (.A(net241),
    .B(_07475_),
    .X(_07477_));
 sky130_fd_sc_hd__nand3_2 _17965_ (.A(_07899_),
    .B(_07459_),
    .C(_07470_),
    .Y(_07478_));
 sky130_fd_sc_hd__o221ai_4 _17966_ (.A1(_07844_),
    .A2(_07866_),
    .B1(_05485_),
    .B2(_07458_),
    .C1(_07474_),
    .Y(_07479_));
 sky130_fd_sc_hd__a21oi_1 _17967_ (.A1(_07044_),
    .A2(_07169_),
    .B1(_07172_),
    .Y(_07480_));
 sky130_fd_sc_hd__a31o_1 _17968_ (.A1(net376),
    .A2(_07022_),
    .A3(_07169_),
    .B1(_07172_),
    .X(_07481_));
 sky130_fd_sc_hd__a32oi_4 _17969_ (.A1(_07167_),
    .A2(_07168_),
    .A3(_07033_),
    .B1(_06849_),
    .B2(_06855_),
    .Y(_07482_));
 sky130_fd_sc_hd__a22oi_2 _17970_ (.A1(_07478_),
    .A2(_07479_),
    .B1(_07481_),
    .B2(_07174_),
    .Y(_07484_));
 sky130_fd_sc_hd__o2bb2ai_1 _17971_ (.A1_N(_07478_),
    .A2_N(_07479_),
    .B1(_07480_),
    .B2(_07173_),
    .Y(_07485_));
 sky130_fd_sc_hd__o21ai_2 _17972_ (.A1(_07175_),
    .A2(_07482_),
    .B1(_07479_),
    .Y(_07486_));
 sky130_fd_sc_hd__o211ai_2 _17973_ (.A1(_07175_),
    .A2(_07482_),
    .B1(_07479_),
    .C1(_07478_),
    .Y(_07487_));
 sky130_fd_sc_hd__o21ai_1 _17974_ (.A1(net266),
    .A2(_05751_),
    .B1(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__nand3_1 _17975_ (.A(_07485_),
    .B(_07487_),
    .C(net241),
    .Y(_07489_));
 sky130_fd_sc_hd__o22ai_4 _17976_ (.A1(net241),
    .A2(_07475_),
    .B1(_07484_),
    .B2(_07488_),
    .Y(_07490_));
 sky130_fd_sc_hd__a211o_2 _17977_ (.A1(_07477_),
    .A2(_07489_),
    .B1(net259),
    .C1(net256),
    .X(_07491_));
 sky130_fd_sc_hd__o32a_1 _17978_ (.A1(net381),
    .A2(_06310_),
    .A3(_07181_),
    .B1(_07189_),
    .B2(_07186_),
    .X(_07492_));
 sky130_fd_sc_hd__o32ai_4 _17979_ (.A1(_06289_),
    .A2(_06310_),
    .A3(_07181_),
    .B1(_07189_),
    .B2(_07186_),
    .Y(_07493_));
 sky130_fd_sc_hd__a31o_1 _17980_ (.A1(_07485_),
    .A2(_07487_),
    .A3(net241),
    .B1(_07044_),
    .X(_07495_));
 sky130_fd_sc_hd__a311oi_1 _17981_ (.A1(_07485_),
    .A2(_07487_),
    .A3(net241),
    .B1(_07476_),
    .C1(_07044_),
    .Y(_07496_));
 sky130_fd_sc_hd__a2bb2oi_2 _17982_ (.A1_N(_06945_),
    .A2_N(_06967_),
    .B1(_07477_),
    .B2(_07489_),
    .Y(_07497_));
 sky130_fd_sc_hd__o21ai_1 _17983_ (.A1(_06945_),
    .A2(_06967_),
    .B1(_07490_),
    .Y(_07498_));
 sky130_fd_sc_hd__o211ai_2 _17984_ (.A1(_07476_),
    .A2(_07495_),
    .B1(_07498_),
    .C1(_07493_),
    .Y(_07499_));
 sky130_fd_sc_hd__o21ai_1 _17985_ (.A1(_07496_),
    .A2(_07497_),
    .B1(_07492_),
    .Y(_07500_));
 sky130_fd_sc_hd__o211ai_4 _17986_ (.A1(net259),
    .A2(net256),
    .B1(_07499_),
    .C1(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__a21oi_1 _17987_ (.A1(_07491_),
    .A2(_07501_),
    .B1(net212),
    .Y(_07502_));
 sky130_fd_sc_hd__a2bb2oi_2 _17988_ (.A1_N(net394),
    .A2_N(_06267_),
    .B1(_07491_),
    .B2(_07501_),
    .Y(_07503_));
 sky130_fd_sc_hd__o211a_1 _17989_ (.A1(net381),
    .A2(_06310_),
    .B1(_07491_),
    .C1(_07501_),
    .X(_07504_));
 sky130_fd_sc_hd__o211ai_2 _17990_ (.A1(net381),
    .A2(_06310_),
    .B1(_07491_),
    .C1(_07501_),
    .Y(_07506_));
 sky130_fd_sc_hd__a21boi_2 _17991_ (.A1(_07194_),
    .A2(_07200_),
    .B1_N(_07199_),
    .Y(_07507_));
 sky130_fd_sc_hd__o21bai_2 _17992_ (.A1(_07503_),
    .A2(_07504_),
    .B1_N(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__and2_1 _17993_ (.A(_07507_),
    .B(_07506_),
    .X(_07509_));
 sky130_fd_sc_hd__nand3b_1 _17994_ (.A_N(_07503_),
    .B(_07506_),
    .C(_07507_),
    .Y(_07510_));
 sky130_fd_sc_hd__a2bb2oi_1 _17995_ (.A1_N(_06291_),
    .A2_N(_06292_),
    .B1(_07508_),
    .B2(_07510_),
    .Y(_07511_));
 sky130_fd_sc_hd__and3_1 _17996_ (.A(_06294_),
    .B(_07491_),
    .C(_07501_),
    .X(_07512_));
 sky130_fd_sc_hd__a31o_2 _17997_ (.A1(_07508_),
    .A2(_07510_),
    .A3(net212),
    .B1(_07502_),
    .X(_07513_));
 sky130_fd_sc_hd__o311a_1 _17998_ (.A1(_05556_),
    .A2(_06886_),
    .A3(_06890_),
    .B1(_07203_),
    .C1(_07205_),
    .X(_07514_));
 sky130_fd_sc_hd__nand3_1 _17999_ (.A(_07203_),
    .B(_07205_),
    .C(_07207_),
    .Y(_07515_));
 sky130_fd_sc_hd__o211ai_4 _18000_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_07210_),
    .C1(_07515_),
    .Y(_07517_));
 sky130_fd_sc_hd__o22a_1 _18001_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_07208_),
    .B2(_07514_),
    .X(_07518_));
 sky130_fd_sc_hd__o22ai_4 _18002_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_07208_),
    .B2(_07514_),
    .Y(_07519_));
 sky130_fd_sc_hd__o211ai_2 _18003_ (.A1(_06608_),
    .A2(net237),
    .B1(_07517_),
    .C1(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__o21a_1 _18004_ (.A1(_07511_),
    .A2(_07512_),
    .B1(_07520_),
    .X(_07521_));
 sky130_fd_sc_hd__o21ai_2 _18005_ (.A1(_07511_),
    .A2(_07512_),
    .B1(_07520_),
    .Y(_07522_));
 sky130_fd_sc_hd__and4_1 _18006_ (.A(_07513_),
    .B(_07517_),
    .C(_07519_),
    .D(_06612_),
    .X(_07523_));
 sky130_fd_sc_hd__nand4_4 _18007_ (.A(_07513_),
    .B(_07517_),
    .C(_07519_),
    .D(_06612_),
    .Y(_07524_));
 sky130_fd_sc_hd__a311oi_2 _18008_ (.A1(_07508_),
    .A2(_07510_),
    .A3(net212),
    .B1(_07502_),
    .C1(_05862_),
    .Y(_07525_));
 sky130_fd_sc_hd__o21ai_2 _18009_ (.A1(_05239_),
    .A2(_07214_),
    .B1(_07222_),
    .Y(_07526_));
 sky130_fd_sc_hd__o22ai_1 _18010_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_07217_),
    .B2(_07221_),
    .Y(_07528_));
 sky130_fd_sc_hd__o211ai_2 _18011_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_07218_),
    .C1(_07222_),
    .Y(_07529_));
 sky130_fd_sc_hd__nand3_2 _18012_ (.A(_07528_),
    .B(_07529_),
    .C(net208),
    .Y(_07530_));
 sky130_fd_sc_hd__o21ai_1 _18013_ (.A1(_07521_),
    .A2(_07523_),
    .B1(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__o2111ai_4 _18014_ (.A1(_03399_),
    .A2(_05491_),
    .B1(net396),
    .C1(_07522_),
    .D1(_07524_),
    .Y(_07532_));
 sky130_fd_sc_hd__o31ai_4 _18015_ (.A1(_07521_),
    .A2(_07523_),
    .A3(_07530_),
    .B1(_07531_),
    .Y(_07533_));
 sky130_fd_sc_hd__a31oi_4 _18016_ (.A1(_07223_),
    .A2(_07224_),
    .A3(net1),
    .B1(_05239_),
    .Y(_07534_));
 sky130_fd_sc_hd__or2_1 _18017_ (.A(_05250_),
    .B(_07235_),
    .X(_07535_));
 sky130_fd_sc_hd__a41o_1 _18018_ (.A1(_07223_),
    .A2(_07224_),
    .A3(net1),
    .A4(_05239_),
    .B1(_07232_),
    .X(_07536_));
 sky130_fd_sc_hd__o21ai_1 _18019_ (.A1(_07534_),
    .A2(_07536_),
    .B1(_07533_),
    .Y(_07537_));
 sky130_fd_sc_hd__o31ai_1 _18020_ (.A1(_07533_),
    .A2(_07534_),
    .A3(_07536_),
    .B1(_07537_),
    .Y(_07539_));
 sky130_fd_sc_hd__o311a_1 _18021_ (.A1(_07533_),
    .A2(_07534_),
    .A3(_07536_),
    .B1(net1),
    .C1(_07537_),
    .X(_07540_));
 sky130_fd_sc_hd__or2_2 _18022_ (.A(_03289_),
    .B(_07539_),
    .X(_07541_));
 sky130_fd_sc_hd__and2_1 _18023_ (.A(_03289_),
    .B(_07539_),
    .X(_07542_));
 sky130_fd_sc_hd__o21ai_4 _18024_ (.A1(net45),
    .A2(_07226_),
    .B1(net409),
    .Y(_07543_));
 sky130_fd_sc_hd__and2_4 _18025_ (.A(_07543_),
    .B(net46),
    .X(_07544_));
 sky130_fd_sc_hd__nand2_8 _18026_ (.A(_07543_),
    .B(net46),
    .Y(_07545_));
 sky130_fd_sc_hd__nor2_8 _18027_ (.A(net46),
    .B(_07543_),
    .Y(_07546_));
 sky130_fd_sc_hd__or2_4 _18028_ (.A(net46),
    .B(_07543_),
    .X(_07547_));
 sky130_fd_sc_hd__nand2_8 _18029_ (.A(_07545_),
    .B(_07547_),
    .Y(_07548_));
 sky130_fd_sc_hd__nor2_8 _18030_ (.A(_07544_),
    .B(net184),
    .Y(_07550_));
 sky130_fd_sc_hd__or3_1 _18031_ (.A(_07544_),
    .B(net184),
    .C(_07539_),
    .X(_07551_));
 sky130_fd_sc_hd__o31a_1 _18032_ (.A1(_07540_),
    .A2(_07550_),
    .A3(_07542_),
    .B1(_07551_),
    .X(_07552_));
 sky130_fd_sc_hd__xnor2_1 _18033_ (.A(_07239_),
    .B(_07552_),
    .Y(net78));
 sky130_fd_sc_hd__nand3_1 _18034_ (.A(_06908_),
    .B(_07236_),
    .C(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__or3_4 _18035_ (.A(net13),
    .B(net14),
    .C(_06913_),
    .X(_07554_));
 sky130_fd_sc_hd__and3b_4 _18036_ (.A_N(net15),
    .B(_07554_),
    .C(net410),
    .X(_07555_));
 sky130_fd_sc_hd__or3b_4 _18037_ (.A(_03399_),
    .B(net15),
    .C_N(_07554_),
    .X(_07556_));
 sky130_fd_sc_hd__a21boi_4 _18038_ (.A1(_07554_),
    .A2(net410),
    .B1_N(net15),
    .Y(_07557_));
 sky130_fd_sc_hd__a21bo_4 _18039_ (.A1(_07554_),
    .A2(net410),
    .B1_N(net15),
    .X(_07558_));
 sky130_fd_sc_hd__o311a_4 _18040_ (.A1(net13),
    .A2(net14),
    .A3(_06913_),
    .B1(net15),
    .C1(net410),
    .X(_07560_));
 sky130_fd_sc_hd__o211ai_4 _18041_ (.A1(net14),
    .A2(_07240_),
    .B1(net15),
    .C1(net410),
    .Y(_07561_));
 sky130_fd_sc_hd__a21oi_4 _18042_ (.A1(_07554_),
    .A2(net410),
    .B1(net15),
    .Y(_07562_));
 sky130_fd_sc_hd__a21o_4 _18043_ (.A1(_07554_),
    .A2(net410),
    .B1(net15),
    .X(_07563_));
 sky130_fd_sc_hd__nand2_8 _18044_ (.A(_07561_),
    .B(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__nor2_8 _18045_ (.A(_07560_),
    .B(net217),
    .Y(_07565_));
 sky130_fd_sc_hd__or3_2 _18046_ (.A(_03178_),
    .B(_07560_),
    .C(_07562_),
    .X(_07566_));
 sky130_fd_sc_hd__a31o_1 _18047_ (.A1(net33),
    .A2(_07561_),
    .A3(_07563_),
    .B1(net222),
    .X(_07567_));
 sky130_fd_sc_hd__o221ai_4 _18048_ (.A1(net234),
    .A2(_06925_),
    .B1(_07249_),
    .B2(net227),
    .C1(_06933_),
    .Y(_07568_));
 sky130_fd_sc_hd__or4_1 _18049_ (.A(_03178_),
    .B(_07244_),
    .C(_07245_),
    .D(_07564_),
    .X(_07569_));
 sky130_fd_sc_hd__o31a_1 _18050_ (.A1(_07560_),
    .A2(_07562_),
    .A3(_07249_),
    .B1(_07567_),
    .X(_07571_));
 sky130_fd_sc_hd__o21ai_2 _18051_ (.A1(_07564_),
    .A2(_07249_),
    .B1(_07567_),
    .Y(_07572_));
 sky130_fd_sc_hd__o211ai_4 _18052_ (.A1(net225),
    .A2(_07248_),
    .B1(_07571_),
    .C1(_07568_),
    .Y(_07573_));
 sky130_fd_sc_hd__o211ai_4 _18053_ (.A1(_07253_),
    .A2(_07254_),
    .B1(_07572_),
    .C1(_07250_),
    .Y(_07574_));
 sky130_fd_sc_hd__o221a_2 _18054_ (.A1(_05130_),
    .A2(_05152_),
    .B1(_07555_),
    .B2(_07557_),
    .C1(net33),
    .X(_07575_));
 sky130_fd_sc_hd__a31o_1 _18055_ (.A1(_07574_),
    .A2(net405),
    .A3(_07573_),
    .B1(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__a31oi_4 _18056_ (.A1(_07574_),
    .A2(net405),
    .A3(_07573_),
    .B1(_07575_),
    .Y(_07577_));
 sky130_fd_sc_hd__or3_2 _18057_ (.A(_05348_),
    .B(net401),
    .C(_07577_),
    .X(_07578_));
 sky130_fd_sc_hd__a21oi_2 _18058_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_07577_),
    .Y(_07579_));
 sky130_fd_sc_hd__o21ai_1 _18059_ (.A1(_06914_),
    .A2(_06916_),
    .B1(_07576_),
    .Y(_07580_));
 sky130_fd_sc_hd__and3_1 _18060_ (.A(_06915_),
    .B(_06917_),
    .C(_07577_),
    .X(_07582_));
 sky130_fd_sc_hd__a311o_1 _18061_ (.A1(_07574_),
    .A2(net405),
    .A3(_07573_),
    .B1(_07575_),
    .C1(net225),
    .X(_07583_));
 sky130_fd_sc_hd__nor2_1 _18062_ (.A(_07579_),
    .B(_07582_),
    .Y(_07584_));
 sky130_fd_sc_hd__nand2_1 _18063_ (.A(_07580_),
    .B(_07583_),
    .Y(_07585_));
 sky130_fd_sc_hd__nand4_4 _18064_ (.A(_06946_),
    .B(_06647_),
    .C(_06341_),
    .D(_06942_),
    .Y(_07586_));
 sky130_fd_sc_hd__o221ai_4 _18065_ (.A1(_06349_),
    .A2(_06352_),
    .B1(_07265_),
    .B2(_07259_),
    .C1(_07264_),
    .Y(_07587_));
 sky130_fd_sc_hd__nor2_2 _18066_ (.A(_07586_),
    .B(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__a211o_1 _18067_ (.A1(_06350_),
    .A2(_06353_),
    .B1(_07267_),
    .C1(_07586_),
    .X(_07589_));
 sky130_fd_sc_hd__o22ai_2 _18068_ (.A1(_07259_),
    .A2(_07265_),
    .B1(_07262_),
    .B2(_07586_),
    .Y(_07590_));
 sky130_fd_sc_hd__a21oi_4 _18069_ (.A1(_07268_),
    .A2(_07266_),
    .B1(_07590_),
    .Y(_07591_));
 sky130_fd_sc_hd__a21o_1 _18070_ (.A1(_07268_),
    .A2(_07266_),
    .B1(_07590_),
    .X(_07593_));
 sky130_fd_sc_hd__o21ai_2 _18071_ (.A1(_07586_),
    .A2(_07587_),
    .B1(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__o22a_1 _18072_ (.A1(_07579_),
    .A2(_07582_),
    .B1(_07588_),
    .B2(_07591_),
    .X(_07595_));
 sky130_fd_sc_hd__o22ai_2 _18073_ (.A1(_07579_),
    .A2(_07582_),
    .B1(_07588_),
    .B2(_07591_),
    .Y(_07596_));
 sky130_fd_sc_hd__nand3_2 _18074_ (.A(_07593_),
    .B(_07584_),
    .C(_07589_),
    .Y(_07597_));
 sky130_fd_sc_hd__o31ai_2 _18075_ (.A1(_07585_),
    .A2(_07588_),
    .A3(_07591_),
    .B1(_05403_),
    .Y(_07598_));
 sky130_fd_sc_hd__nand3_2 _18076_ (.A(_05403_),
    .B(_07596_),
    .C(_07597_),
    .Y(_07599_));
 sky130_fd_sc_hd__o22ai_4 _18077_ (.A1(_05403_),
    .A2(_07577_),
    .B1(_07595_),
    .B2(_07598_),
    .Y(_07600_));
 sky130_fd_sc_hd__a2bb2oi_2 _18078_ (.A1_N(_06622_),
    .A2_N(_06624_),
    .B1(_07578_),
    .B2(_07599_),
    .Y(_07601_));
 sky130_fd_sc_hd__o21ai_4 _18079_ (.A1(_06622_),
    .A2(_06624_),
    .B1(_07600_),
    .Y(_07602_));
 sky130_fd_sc_hd__a31oi_1 _18080_ (.A1(_05403_),
    .A2(_07596_),
    .A3(_07597_),
    .B1(net232),
    .Y(_07604_));
 sky130_fd_sc_hd__o211a_1 _18081_ (.A1(_05403_),
    .A2(_07577_),
    .B1(net234),
    .C1(_07599_),
    .X(_07605_));
 sky130_fd_sc_hd__o211ai_4 _18082_ (.A1(_05403_),
    .A2(_07577_),
    .B1(net234),
    .C1(_07599_),
    .Y(_07606_));
 sky130_fd_sc_hd__a21oi_2 _18083_ (.A1(_07578_),
    .A2(_07604_),
    .B1(_07601_),
    .Y(_07607_));
 sky130_fd_sc_hd__o221ai_4 _18084_ (.A1(_06314_),
    .A2(_07275_),
    .B1(_06959_),
    .B2(_06960_),
    .C1(_06955_),
    .Y(_07608_));
 sky130_fd_sc_hd__o21ai_2 _18085_ (.A1(net251),
    .A2(_07276_),
    .B1(_07608_),
    .Y(_07609_));
 sky130_fd_sc_hd__nand4b_4 _18086_ (.A_N(_07279_),
    .B(_07602_),
    .C(_07606_),
    .D(_07608_),
    .Y(_07610_));
 sky130_fd_sc_hd__o21ai_4 _18087_ (.A1(_07601_),
    .A2(_07605_),
    .B1(_07609_),
    .Y(_07611_));
 sky130_fd_sc_hd__nand3_2 _18088_ (.A(_07611_),
    .B(net359),
    .C(_07610_),
    .Y(_07612_));
 sky130_fd_sc_hd__and3_2 _18089_ (.A(_05687_),
    .B(_05709_),
    .C(_07600_),
    .X(_07613_));
 sky130_fd_sc_hd__a211o_2 _18090_ (.A1(_07578_),
    .A2(_07599_),
    .B1(_05676_),
    .C1(_05698_),
    .X(_07615_));
 sky130_fd_sc_hd__a31o_1 _18091_ (.A1(_07610_),
    .A2(_07611_),
    .A3(net359),
    .B1(_07613_),
    .X(_07616_));
 sky130_fd_sc_hd__a21oi_4 _18092_ (.A1(_07612_),
    .A2(_07615_),
    .B1(_06314_),
    .Y(_07617_));
 sky130_fd_sc_hd__a22o_1 _18093_ (.A1(_06306_),
    .A2(_06308_),
    .B1(_07612_),
    .B2(_07615_),
    .X(_07618_));
 sky130_fd_sc_hd__a31oi_1 _18094_ (.A1(_07610_),
    .A2(_07611_),
    .A3(net359),
    .B1(net251),
    .Y(_07619_));
 sky130_fd_sc_hd__a31o_1 _18095_ (.A1(_07610_),
    .A2(_07611_),
    .A3(net359),
    .B1(net251),
    .X(_07620_));
 sky130_fd_sc_hd__a311oi_4 _18096_ (.A1(_07610_),
    .A2(_07611_),
    .A3(net359),
    .B1(_07613_),
    .C1(net251),
    .Y(_07621_));
 sky130_fd_sc_hd__a311o_1 _18097_ (.A1(_07610_),
    .A2(_07611_),
    .A3(net359),
    .B1(_07613_),
    .C1(net251),
    .X(_07622_));
 sky130_fd_sc_hd__a21oi_2 _18098_ (.A1(_07615_),
    .A2(_07619_),
    .B1(_07617_),
    .Y(_07623_));
 sky130_fd_sc_hd__o21ai_1 _18099_ (.A1(_07613_),
    .A2(_07620_),
    .B1(_07618_),
    .Y(_07624_));
 sky130_fd_sc_hd__o22ai_2 _18100_ (.A1(net254),
    .A2(_07290_),
    .B1(_07299_),
    .B2(_07301_),
    .Y(_07626_));
 sky130_fd_sc_hd__o221a_1 _18101_ (.A1(net254),
    .A2(_07290_),
    .B1(_07617_),
    .B2(_07621_),
    .C1(_07302_),
    .X(_07627_));
 sky130_fd_sc_hd__o221ai_4 _18102_ (.A1(_07290_),
    .A2(net254),
    .B1(_07621_),
    .B2(_07617_),
    .C1(_07302_),
    .Y(_07628_));
 sky130_fd_sc_hd__a21oi_1 _18103_ (.A1(_07293_),
    .A2(_07302_),
    .B1(_07624_),
    .Y(_07629_));
 sky130_fd_sc_hd__nand2_1 _18104_ (.A(_07626_),
    .B(_07623_),
    .Y(_07630_));
 sky130_fd_sc_hd__o21ai_2 _18105_ (.A1(_07627_),
    .A2(_07629_),
    .B1(net357),
    .Y(_07631_));
 sky130_fd_sc_hd__a211o_2 _18106_ (.A1(_07612_),
    .A2(_07615_),
    .B1(net379),
    .C1(net378),
    .X(_07632_));
 sky130_fd_sc_hd__inv_2 _18107_ (.A(_07632_),
    .Y(_07633_));
 sky130_fd_sc_hd__nand3_2 _18108_ (.A(_07630_),
    .B(net357),
    .C(_07628_),
    .Y(_07634_));
 sky130_fd_sc_hd__a2bb2oi_2 _18109_ (.A1_N(_06009_),
    .A2_N(_06010_),
    .B1(_07632_),
    .B2(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__o211ai_4 _18110_ (.A1(_07616_),
    .A2(net357),
    .B1(net253),
    .C1(_07631_),
    .Y(_07637_));
 sky130_fd_sc_hd__a311oi_4 _18111_ (.A1(_07630_),
    .A2(net357),
    .A3(_07628_),
    .B1(_07633_),
    .C1(net253),
    .Y(_07638_));
 sky130_fd_sc_hd__o211ai_4 _18112_ (.A1(net286),
    .A2(_06012_),
    .B1(_07632_),
    .C1(_07634_),
    .Y(_07639_));
 sky130_fd_sc_hd__o21ai_2 _18113_ (.A1(_07309_),
    .A2(_07313_),
    .B1(_07308_),
    .Y(_07640_));
 sky130_fd_sc_hd__a21oi_2 _18114_ (.A1(_07312_),
    .A2(_07310_),
    .B1(_07306_),
    .Y(_07641_));
 sky130_fd_sc_hd__o21ai_4 _18115_ (.A1(_07635_),
    .A2(_07638_),
    .B1(_07641_),
    .Y(_07642_));
 sky130_fd_sc_hd__nand3_4 _18116_ (.A(_07640_),
    .B(_07639_),
    .C(_07637_),
    .Y(_07643_));
 sky130_fd_sc_hd__o311a_2 _18117_ (.A1(_06793_),
    .A2(_07616_),
    .A3(_06815_),
    .B1(_07724_),
    .C1(_07631_),
    .X(_07644_));
 sky130_fd_sc_hd__a211o_1 _18118_ (.A1(_07632_),
    .A2(_07634_),
    .B1(net373),
    .C1(net371),
    .X(_07645_));
 sky130_fd_sc_hd__o211ai_2 _18119_ (.A1(net373),
    .A2(net371),
    .B1(_07642_),
    .C1(_07643_),
    .Y(_07646_));
 sky130_fd_sc_hd__a31o_1 _18120_ (.A1(_07642_),
    .A2(_07643_),
    .A3(net355),
    .B1(_07644_),
    .X(_07648_));
 sky130_fd_sc_hd__a31oi_2 _18121_ (.A1(_07642_),
    .A2(_07643_),
    .A3(net355),
    .B1(_07644_),
    .Y(_07649_));
 sky130_fd_sc_hd__a311o_1 _18122_ (.A1(_07642_),
    .A2(_07643_),
    .A3(net355),
    .B1(_07644_),
    .C1(net338),
    .X(_07650_));
 sky130_fd_sc_hd__a311oi_4 _18123_ (.A1(_07642_),
    .A2(_07643_),
    .A3(net355),
    .B1(_07644_),
    .C1(net261),
    .Y(_07651_));
 sky130_fd_sc_hd__a311o_1 _18124_ (.A1(_07642_),
    .A2(_07643_),
    .A3(net355),
    .B1(_07644_),
    .C1(net261),
    .X(_07652_));
 sky130_fd_sc_hd__a2bb2oi_2 _18125_ (.A1_N(_05760_),
    .A2_N(net290),
    .B1(_07645_),
    .B2(_07646_),
    .Y(_07653_));
 sky130_fd_sc_hd__o21ai_4 _18126_ (.A1(_05760_),
    .A2(net290),
    .B1(_07648_),
    .Y(_07654_));
 sky130_fd_sc_hd__nor2_1 _18127_ (.A(_07651_),
    .B(_07653_),
    .Y(_07655_));
 sky130_fd_sc_hd__and3_1 _18128_ (.A(_06415_),
    .B(_06709_),
    .C(_06710_),
    .X(_07656_));
 sky130_fd_sc_hd__nand4b_2 _18129_ (.A_N(_06427_),
    .B(_07020_),
    .C(_07025_),
    .D(_07656_),
    .Y(_07657_));
 sky130_fd_sc_hd__nand3_1 _18130_ (.A(_07026_),
    .B(_07326_),
    .C(_07656_),
    .Y(_07659_));
 sky130_fd_sc_hd__nor2_1 _18131_ (.A(_07328_),
    .B(_07657_),
    .Y(_07660_));
 sky130_fd_sc_hd__nand3b_2 _18132_ (.A_N(_07657_),
    .B(_07327_),
    .C(_07326_),
    .Y(_07661_));
 sky130_fd_sc_hd__o211a_2 _18133_ (.A1(_07331_),
    .A2(_07325_),
    .B1(_07327_),
    .C1(_07659_),
    .X(_07662_));
 sky130_fd_sc_hd__o211ai_2 _18134_ (.A1(_07331_),
    .A2(_07325_),
    .B1(_07327_),
    .C1(_07659_),
    .Y(_07663_));
 sky130_fd_sc_hd__a31o_1 _18135_ (.A1(_07327_),
    .A2(_07335_),
    .A3(_07659_),
    .B1(_07660_),
    .X(_07664_));
 sky130_fd_sc_hd__nand4_4 _18136_ (.A(_07652_),
    .B(_07654_),
    .C(_07661_),
    .D(_07663_),
    .Y(_07665_));
 sky130_fd_sc_hd__o22ai_4 _18137_ (.A1(_07651_),
    .A2(_07653_),
    .B1(_07660_),
    .B2(_07662_),
    .Y(_07666_));
 sky130_fd_sc_hd__o21ai_1 _18138_ (.A1(_07660_),
    .A2(_07662_),
    .B1(_07655_),
    .Y(_07667_));
 sky130_fd_sc_hd__o211ai_1 _18139_ (.A1(_07651_),
    .A2(_07653_),
    .B1(_07661_),
    .C1(_07663_),
    .Y(_07668_));
 sky130_fd_sc_hd__nand3_2 _18140_ (.A(_07667_),
    .B(_07668_),
    .C(net338),
    .Y(_07670_));
 sky130_fd_sc_hd__a21o_2 _18141_ (.A1(_07645_),
    .A2(_07646_),
    .B1(net338),
    .X(_07671_));
 sky130_fd_sc_hd__inv_2 _18142_ (.A(_07671_),
    .Y(_07672_));
 sky130_fd_sc_hd__nand3_2 _18143_ (.A(_07666_),
    .B(net338),
    .C(_07665_),
    .Y(_07673_));
 sky130_fd_sc_hd__and3_2 _18144_ (.A(_09840_),
    .B(_07650_),
    .C(_07670_),
    .X(_07674_));
 sky130_fd_sc_hd__a211o_1 _18145_ (.A1(_07671_),
    .A2(_07673_),
    .B1(_09785_),
    .C1(net349),
    .X(_07675_));
 sky130_fd_sc_hd__a311oi_4 _18146_ (.A1(_07666_),
    .A2(net338),
    .A3(_07665_),
    .B1(_07672_),
    .C1(net291),
    .Y(_07676_));
 sky130_fd_sc_hd__nand3_4 _18147_ (.A(_07673_),
    .B(net267),
    .C(_07671_),
    .Y(_07677_));
 sky130_fd_sc_hd__a2bb2oi_1 _18148_ (.A1_N(_05500_),
    .A2_N(_05503_),
    .B1(_07671_),
    .B2(_07673_),
    .Y(_07678_));
 sky130_fd_sc_hd__o211ai_4 _18149_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_07650_),
    .C1(_07670_),
    .Y(_07679_));
 sky130_fd_sc_hd__o211a_1 _18150_ (.A1(_07046_),
    .A2(_07042_),
    .B1(_07041_),
    .C1(_07346_),
    .X(_07681_));
 sky130_fd_sc_hd__o21ai_1 _18151_ (.A1(_07343_),
    .A2(_07342_),
    .B1(_07346_),
    .Y(_07682_));
 sky130_fd_sc_hd__a21oi_2 _18152_ (.A1(_07341_),
    .A2(_07344_),
    .B1(_07345_),
    .Y(_07683_));
 sky130_fd_sc_hd__o2bb2ai_2 _18153_ (.A1_N(_07677_),
    .A2_N(_07679_),
    .B1(_07681_),
    .B2(_07343_),
    .Y(_07684_));
 sky130_fd_sc_hd__nand3_2 _18154_ (.A(_07677_),
    .B(_07679_),
    .C(_07682_),
    .Y(_07685_));
 sky130_fd_sc_hd__o311a_1 _18155_ (.A1(_07683_),
    .A2(_07678_),
    .A3(_07676_),
    .B1(net336),
    .C1(_07684_),
    .X(_07686_));
 sky130_fd_sc_hd__nand3_1 _18156_ (.A(_07684_),
    .B(_07685_),
    .C(net336),
    .Y(_07687_));
 sky130_fd_sc_hd__nor2_1 _18157_ (.A(_07674_),
    .B(_07686_),
    .Y(_07688_));
 sky130_fd_sc_hd__inv_2 _18158_ (.A(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__o221a_1 _18159_ (.A1(_02137_),
    .A2(_07056_),
    .B1(_07068_),
    .B2(_07079_),
    .C1(_07359_),
    .X(_07690_));
 sky130_fd_sc_hd__a21oi_1 _18160_ (.A1(_07059_),
    .A2(_07080_),
    .B1(_07361_),
    .Y(_07692_));
 sky130_fd_sc_hd__o21ai_1 _18161_ (.A1(_07361_),
    .A2(_07365_),
    .B1(_07359_),
    .Y(_07693_));
 sky130_fd_sc_hd__a31oi_1 _18162_ (.A1(_07684_),
    .A2(_07685_),
    .A3(net336),
    .B1(net293),
    .Y(_07694_));
 sky130_fd_sc_hd__a311oi_2 _18163_ (.A1(_07684_),
    .A2(_07685_),
    .A3(net336),
    .B1(net293),
    .C1(_07674_),
    .Y(_07695_));
 sky130_fd_sc_hd__a311o_2 _18164_ (.A1(_07684_),
    .A2(_07685_),
    .A3(net336),
    .B1(net293),
    .C1(_07674_),
    .X(_07696_));
 sky130_fd_sc_hd__a2bb2oi_2 _18165_ (.A1_N(_05242_),
    .A2_N(net314),
    .B1(_07675_),
    .B2(_07687_),
    .Y(_07697_));
 sky130_fd_sc_hd__o22ai_2 _18166_ (.A1(_05242_),
    .A2(net314),
    .B1(_07674_),
    .B2(_07686_),
    .Y(_07698_));
 sky130_fd_sc_hd__o211ai_1 _18167_ (.A1(_07361_),
    .A2(_07690_),
    .B1(_07696_),
    .C1(_07698_),
    .Y(_07699_));
 sky130_fd_sc_hd__o22ai_1 _18168_ (.A1(_07358_),
    .A2(_07692_),
    .B1(_07695_),
    .B2(_07697_),
    .Y(_07700_));
 sky130_fd_sc_hd__o211ai_1 _18169_ (.A1(_07358_),
    .A2(_07692_),
    .B1(_07696_),
    .C1(_07698_),
    .Y(_07701_));
 sky130_fd_sc_hd__o22ai_1 _18170_ (.A1(_07361_),
    .A2(_07690_),
    .B1(_07695_),
    .B2(_07697_),
    .Y(_07703_));
 sky130_fd_sc_hd__nand3_2 _18171_ (.A(_07699_),
    .B(_07700_),
    .C(net334),
    .Y(_07704_));
 sky130_fd_sc_hd__a211o_1 _18172_ (.A1(_07675_),
    .A2(_07687_),
    .B1(net347),
    .C1(net346),
    .X(_07705_));
 sky130_fd_sc_hd__nand3_2 _18173_ (.A(_07701_),
    .B(_07703_),
    .C(net334),
    .Y(_07706_));
 sky130_fd_sc_hd__o21ai_1 _18174_ (.A1(net333),
    .A2(_07688_),
    .B1(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__and3_1 _18175_ (.A(_07706_),
    .B(net299),
    .C(_07705_),
    .X(_07708_));
 sky130_fd_sc_hd__nand3_2 _18176_ (.A(_07706_),
    .B(net299),
    .C(_07705_),
    .Y(_07709_));
 sky130_fd_sc_hd__o311a_2 _18177_ (.A1(net334),
    .A2(_07674_),
    .A3(_07686_),
    .B1(_07704_),
    .C1(net298),
    .X(_07710_));
 sky130_fd_sc_hd__o211ai_4 _18178_ (.A1(_07689_),
    .A2(net334),
    .B1(net298),
    .C1(_07704_),
    .Y(_07711_));
 sky130_fd_sc_hd__a22oi_2 _18179_ (.A1(_02148_),
    .A2(_07374_),
    .B1(_07376_),
    .B2(_07090_),
    .Y(_07712_));
 sky130_fd_sc_hd__o32a_1 _18180_ (.A1(_02049_),
    .A2(net342),
    .A3(_07374_),
    .B1(_07377_),
    .B2(_07379_),
    .X(_07714_));
 sky130_fd_sc_hd__o2bb2ai_1 _18181_ (.A1_N(_07709_),
    .A2_N(_07711_),
    .B1(_07712_),
    .B2(_07381_),
    .Y(_07715_));
 sky130_fd_sc_hd__o2111ai_4 _18182_ (.A1(_07377_),
    .A2(_07379_),
    .B1(_07382_),
    .C1(_07709_),
    .D1(_07711_),
    .Y(_07716_));
 sky130_fd_sc_hd__nand3_4 _18183_ (.A(_07715_),
    .B(_07716_),
    .C(net312),
    .Y(_07717_));
 sky130_fd_sc_hd__a211o_2 _18184_ (.A1(_07705_),
    .A2(_07706_),
    .B1(_12670_),
    .C1(_12681_),
    .X(_07718_));
 sky130_fd_sc_hd__nand2_2 _18185_ (.A(_07717_),
    .B(_07718_),
    .Y(_07719_));
 sky130_fd_sc_hd__inv_2 _18186_ (.A(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__a21oi_1 _18187_ (.A1(_07717_),
    .A2(_07718_),
    .B1(_02137_),
    .Y(_07721_));
 sky130_fd_sc_hd__a21o_1 _18188_ (.A1(_07717_),
    .A2(_07718_),
    .B1(_02137_),
    .X(_07722_));
 sky130_fd_sc_hd__and3_1 _18189_ (.A(_07717_),
    .B(_07718_),
    .C(_02137_),
    .X(_07723_));
 sky130_fd_sc_hd__o211ai_2 _18190_ (.A1(_02093_),
    .A2(_02115_),
    .B1(_07717_),
    .C1(_07718_),
    .Y(_07725_));
 sky130_fd_sc_hd__and4_1 _18191_ (.A(_06496_),
    .B(_06499_),
    .C(_06774_),
    .D(_06776_),
    .X(_07726_));
 sky130_fd_sc_hd__nand4_1 _18192_ (.A(_06496_),
    .B(_06499_),
    .C(_06774_),
    .D(_06776_),
    .Y(_07727_));
 sky130_fd_sc_hd__a21oi_1 _18193_ (.A1(net325),
    .A2(_07103_),
    .B1(_07727_),
    .Y(_07728_));
 sky130_fd_sc_hd__nor3_1 _18194_ (.A(_07107_),
    .B(_07727_),
    .C(_07109_),
    .Y(_07729_));
 sky130_fd_sc_hd__nand3_2 _18195_ (.A(_07728_),
    .B(_07396_),
    .C(_07108_),
    .Y(_07730_));
 sky130_fd_sc_hd__o211a_1 _18196_ (.A1(_07401_),
    .A2(_07394_),
    .B1(_07398_),
    .C1(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__o211ai_4 _18197_ (.A1(_07401_),
    .A2(_07394_),
    .B1(_07398_),
    .C1(_07730_),
    .Y(_07732_));
 sky130_fd_sc_hd__nand4_1 _18198_ (.A(_07108_),
    .B(_07111_),
    .C(_07726_),
    .D(_06501_),
    .Y(_07733_));
 sky130_fd_sc_hd__nand4_4 _18199_ (.A(_07396_),
    .B(_07729_),
    .C(_07398_),
    .D(_06501_),
    .Y(_07734_));
 sky130_fd_sc_hd__a41o_1 _18200_ (.A1(_06501_),
    .A2(_07396_),
    .A3(_07398_),
    .A4(_07729_),
    .B1(_07731_),
    .X(_07736_));
 sky130_fd_sc_hd__o31ai_2 _18201_ (.A1(_07394_),
    .A2(_07397_),
    .A3(_07733_),
    .B1(_07725_),
    .Y(_07737_));
 sky130_fd_sc_hd__o2111ai_4 _18202_ (.A1(_02148_),
    .A2(_07719_),
    .B1(_07722_),
    .C1(_07732_),
    .D1(_07734_),
    .Y(_07738_));
 sky130_fd_sc_hd__nor2_1 _18203_ (.A(_07721_),
    .B(_07723_),
    .Y(_07739_));
 sky130_fd_sc_hd__a22o_2 _18204_ (.A1(_07722_),
    .A2(_07725_),
    .B1(_07732_),
    .B2(_07734_),
    .X(_07740_));
 sky130_fd_sc_hd__nand3_2 _18205_ (.A(_07740_),
    .B(net309),
    .C(_07738_),
    .Y(_07741_));
 sky130_fd_sc_hd__and3_4 _18206_ (.A(_00022_),
    .B(_00044_),
    .C(_07719_),
    .X(_07742_));
 sky130_fd_sc_hd__a211o_2 _18207_ (.A1(_07717_),
    .A2(_07718_),
    .B1(net324),
    .C1(_00033_),
    .X(_07743_));
 sky130_fd_sc_hd__a31oi_4 _18208_ (.A1(_07740_),
    .A2(net309),
    .A3(_07738_),
    .B1(_07742_),
    .Y(_07744_));
 sky130_fd_sc_hd__a21oi_2 _18209_ (.A1(_07741_),
    .A2(_07743_),
    .B1(net280),
    .Y(_07745_));
 sky130_fd_sc_hd__or3_2 _18210_ (.A(net306),
    .B(net303),
    .C(_07744_),
    .X(_07747_));
 sky130_fd_sc_hd__a31o_2 _18211_ (.A1(_07740_),
    .A2(net309),
    .A3(_07738_),
    .B1(net319),
    .X(_07748_));
 sky130_fd_sc_hd__a311oi_4 _18212_ (.A1(_07740_),
    .A2(net309),
    .A3(_07738_),
    .B1(_07742_),
    .C1(net319),
    .Y(_07749_));
 sky130_fd_sc_hd__a22oi_4 _18213_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_07741_),
    .B2(_07743_),
    .Y(_07750_));
 sky130_fd_sc_hd__a21o_1 _18214_ (.A1(_07741_),
    .A2(_07743_),
    .B1(net320),
    .X(_07751_));
 sky130_fd_sc_hd__o31ai_4 _18215_ (.A1(_07124_),
    .A2(_07408_),
    .A3(_07409_),
    .B1(_07412_),
    .Y(_07752_));
 sky130_fd_sc_hd__a31o_1 _18216_ (.A1(_07123_),
    .A2(_07129_),
    .A3(_07412_),
    .B1(_07409_),
    .X(_07753_));
 sky130_fd_sc_hd__o21a_1 _18217_ (.A1(_07749_),
    .A2(_07750_),
    .B1(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__o21ai_4 _18218_ (.A1(_07749_),
    .A2(_07750_),
    .B1(_07753_),
    .Y(_07755_));
 sky130_fd_sc_hd__o21ai_2 _18219_ (.A1(net320),
    .A2(_07744_),
    .B1(_07752_),
    .Y(_07756_));
 sky130_fd_sc_hd__o211ai_4 _18220_ (.A1(_07742_),
    .A2(_07748_),
    .B1(_07752_),
    .C1(_07751_),
    .Y(_07757_));
 sky130_fd_sc_hd__o22ai_2 _18221_ (.A1(net306),
    .A2(net303),
    .B1(_07749_),
    .B2(_07756_),
    .Y(_07758_));
 sky130_fd_sc_hd__o211ai_4 _18222_ (.A1(_07749_),
    .A2(_07756_),
    .B1(net280),
    .C1(_07755_),
    .Y(_07759_));
 sky130_fd_sc_hd__o22ai_4 _18223_ (.A1(net280),
    .A2(_07744_),
    .B1(_07754_),
    .B2(_07758_),
    .Y(_07760_));
 sky130_fd_sc_hd__a311o_2 _18224_ (.A1(_07755_),
    .A2(_07757_),
    .A3(net280),
    .B1(net276),
    .C1(_07745_),
    .X(_07761_));
 sky130_fd_sc_hd__o211a_1 _18225_ (.A1(_07137_),
    .A2(_07139_),
    .B1(_07422_),
    .C1(_07136_),
    .X(_07762_));
 sky130_fd_sc_hd__o21ai_1 _18226_ (.A1(_07429_),
    .A2(_07424_),
    .B1(_07422_),
    .Y(_07763_));
 sky130_fd_sc_hd__a31oi_2 _18227_ (.A1(_07755_),
    .A2(_07757_),
    .A3(net280),
    .B1(net325),
    .Y(_07764_));
 sky130_fd_sc_hd__a311oi_4 _18228_ (.A1(_07755_),
    .A2(_07757_),
    .A3(net280),
    .B1(_07745_),
    .C1(net325),
    .Y(_07765_));
 sky130_fd_sc_hd__o221ai_4 _18229_ (.A1(_12867_),
    .A2(_12877_),
    .B1(net280),
    .B2(_07744_),
    .C1(_07759_),
    .Y(_07766_));
 sky130_fd_sc_hd__a2bb2oi_4 _18230_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_07747_),
    .B2(_07759_),
    .Y(_07768_));
 sky130_fd_sc_hd__o21ai_1 _18231_ (.A1(_12845_),
    .A2(_12856_),
    .B1(_07760_),
    .Y(_07769_));
 sky130_fd_sc_hd__a21oi_1 _18232_ (.A1(_07747_),
    .A2(_07764_),
    .B1(_07768_),
    .Y(_07770_));
 sky130_fd_sc_hd__o211ai_2 _18233_ (.A1(_07424_),
    .A2(_07762_),
    .B1(_07766_),
    .C1(_07769_),
    .Y(_07771_));
 sky130_fd_sc_hd__o22ai_2 _18234_ (.A1(_07423_),
    .A2(_07436_),
    .B1(_07765_),
    .B2(_07768_),
    .Y(_07772_));
 sky130_fd_sc_hd__nand3_1 _18235_ (.A(_07769_),
    .B(_07763_),
    .C(_07766_),
    .Y(_07773_));
 sky130_fd_sc_hd__o22ai_1 _18236_ (.A1(_07424_),
    .A2(_07762_),
    .B1(_07765_),
    .B2(_07768_),
    .Y(_07774_));
 sky130_fd_sc_hd__o211ai_4 _18237_ (.A1(net301),
    .A2(net300),
    .B1(_07771_),
    .C1(_07772_),
    .Y(_07775_));
 sky130_fd_sc_hd__a211o_1 _18238_ (.A1(_07747_),
    .A2(_07759_),
    .B1(_04008_),
    .C1(net300),
    .X(_07776_));
 sky130_fd_sc_hd__o211ai_2 _18239_ (.A1(net301),
    .A2(net300),
    .B1(_07773_),
    .C1(_07774_),
    .Y(_07777_));
 sky130_fd_sc_hd__and3_2 _18240_ (.A(_07777_),
    .B(net331),
    .C(_07776_),
    .X(_07779_));
 sky130_fd_sc_hd__nand3_2 _18241_ (.A(_07777_),
    .B(net331),
    .C(_07776_),
    .Y(_07780_));
 sky130_fd_sc_hd__and3_1 _18242_ (.A(net330),
    .B(_07761_),
    .C(_07775_),
    .X(_07781_));
 sky130_fd_sc_hd__o211ai_4 _18243_ (.A1(_07760_),
    .A2(net275),
    .B1(net330),
    .C1(_07775_),
    .Y(_07782_));
 sky130_fd_sc_hd__o31a_1 _18244_ (.A1(_09971_),
    .A2(_09993_),
    .A3(_07440_),
    .B1(_07447_),
    .X(_07783_));
 sky130_fd_sc_hd__o21ai_2 _18245_ (.A1(_07444_),
    .A2(_07447_),
    .B1(_07443_),
    .Y(_07784_));
 sky130_fd_sc_hd__o2bb2ai_4 _18246_ (.A1_N(_07780_),
    .A2_N(_07782_),
    .B1(_07783_),
    .B2(_07444_),
    .Y(_07785_));
 sky130_fd_sc_hd__o211ai_4 _18247_ (.A1(_07442_),
    .A2(_07449_),
    .B1(_07780_),
    .C1(_07782_),
    .Y(_07786_));
 sky130_fd_sc_hd__nand3_2 _18248_ (.A(_07785_),
    .B(_07786_),
    .C(_05233_),
    .Y(_07787_));
 sky130_fd_sc_hd__and3_2 _18249_ (.A(_05234_),
    .B(_07761_),
    .C(_07775_),
    .X(_07788_));
 sky130_fd_sc_hd__a211o_1 _18250_ (.A1(_07776_),
    .A2(_07777_),
    .B1(net297),
    .C1(_05232_),
    .X(_07790_));
 sky130_fd_sc_hd__a31oi_4 _18251_ (.A1(_07785_),
    .A2(_07786_),
    .A3(_05233_),
    .B1(_07788_),
    .Y(_07791_));
 sky130_fd_sc_hd__a31o_2 _18252_ (.A1(_07785_),
    .A2(_07786_),
    .A3(_05233_),
    .B1(_07788_),
    .X(_07792_));
 sky130_fd_sc_hd__and3_1 _18253_ (.A(_05486_),
    .B(_07787_),
    .C(_07790_),
    .X(_07793_));
 sky130_fd_sc_hd__a22oi_4 _18254_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_07787_),
    .B2(_07790_),
    .Y(_07794_));
 sky130_fd_sc_hd__a22o_2 _18255_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_07787_),
    .B2(_07790_),
    .X(_07795_));
 sky130_fd_sc_hd__a311oi_4 _18256_ (.A1(_07785_),
    .A2(_07786_),
    .A3(_05233_),
    .B1(_07788_),
    .C1(net348),
    .Y(_07796_));
 sky130_fd_sc_hd__a311o_2 _18257_ (.A1(_07785_),
    .A2(_07786_),
    .A3(_05233_),
    .B1(_07788_),
    .C1(net348),
    .X(_07797_));
 sky130_fd_sc_hd__a21oi_4 _18258_ (.A1(_07463_),
    .A2(_07465_),
    .B1(_07466_),
    .Y(_07798_));
 sky130_fd_sc_hd__a32o_2 _18259_ (.A1(_08918_),
    .A2(_07441_),
    .A3(_07454_),
    .B1(_07463_),
    .B2(_07465_),
    .X(_07799_));
 sky130_fd_sc_hd__o21ai_4 _18260_ (.A1(_07794_),
    .A2(_07796_),
    .B1(_07799_),
    .Y(_07801_));
 sky130_fd_sc_hd__nand3_2 _18261_ (.A(_07795_),
    .B(_07797_),
    .C(_07798_),
    .Y(_07802_));
 sky130_fd_sc_hd__o211ai_2 _18262_ (.A1(_05481_),
    .A2(net269),
    .B1(_07801_),
    .C1(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__and3_1 _18263_ (.A(_05482_),
    .B(_05484_),
    .C(_07792_),
    .X(_07804_));
 sky130_fd_sc_hd__o21ai_2 _18264_ (.A1(_07794_),
    .A2(_07796_),
    .B1(_07798_),
    .Y(_07805_));
 sky130_fd_sc_hd__a21oi_1 _18265_ (.A1(_10015_),
    .A2(_07791_),
    .B1(_07798_),
    .Y(_07806_));
 sky130_fd_sc_hd__nand3_2 _18266_ (.A(_07795_),
    .B(_07797_),
    .C(_07799_),
    .Y(_07807_));
 sky130_fd_sc_hd__o211ai_2 _18267_ (.A1(_05481_),
    .A2(net269),
    .B1(_07805_),
    .C1(_07807_),
    .Y(_07808_));
 sky130_fd_sc_hd__a31o_1 _18268_ (.A1(_07801_),
    .A2(_07802_),
    .A3(_05485_),
    .B1(_07793_),
    .X(_07809_));
 sky130_fd_sc_hd__o311a_2 _18269_ (.A1(_05481_),
    .A2(_07792_),
    .A3(net269),
    .B1(_05754_),
    .C1(_07803_),
    .X(_07810_));
 sky130_fd_sc_hd__a311o_1 _18270_ (.A1(_07801_),
    .A2(_07802_),
    .A3(_05485_),
    .B1(net241),
    .C1(_07793_),
    .X(_07812_));
 sky130_fd_sc_hd__o21ai_4 _18271_ (.A1(_07888_),
    .A2(_07475_),
    .B1(_07486_),
    .Y(_07813_));
 sky130_fd_sc_hd__a311oi_4 _18272_ (.A1(_07805_),
    .A2(_07807_),
    .A3(_05485_),
    .B1(_07804_),
    .C1(_08918_),
    .Y(_07814_));
 sky130_fd_sc_hd__o211ai_4 _18273_ (.A1(_05485_),
    .A2(_07791_),
    .B1(_08907_),
    .C1(_07808_),
    .Y(_07815_));
 sky130_fd_sc_hd__a311oi_4 _18274_ (.A1(_07801_),
    .A2(_07802_),
    .A3(_05485_),
    .B1(_07793_),
    .C1(_08907_),
    .Y(_07816_));
 sky130_fd_sc_hd__o211ai_2 _18275_ (.A1(_07792_),
    .A2(_05485_),
    .B1(_08918_),
    .C1(_07803_),
    .Y(_07817_));
 sky130_fd_sc_hd__o2111ai_1 _18276_ (.A1(_07888_),
    .A2(_07475_),
    .B1(_07486_),
    .C1(_07815_),
    .D1(_07817_),
    .Y(_07818_));
 sky130_fd_sc_hd__o21ai_1 _18277_ (.A1(_07814_),
    .A2(_07816_),
    .B1(_07813_),
    .Y(_07819_));
 sky130_fd_sc_hd__nand3_4 _18278_ (.A(_07813_),
    .B(_07815_),
    .C(_07817_),
    .Y(_07820_));
 sky130_fd_sc_hd__o21bai_4 _18279_ (.A1(_07814_),
    .A2(_07816_),
    .B1_N(_07813_),
    .Y(_07821_));
 sky130_fd_sc_hd__a2bb2oi_1 _18280_ (.A1_N(net266),
    .A2_N(_05751_),
    .B1(_07818_),
    .B2(_07819_),
    .Y(_07823_));
 sky130_fd_sc_hd__o211ai_4 _18281_ (.A1(net266),
    .A2(_05751_),
    .B1(_07820_),
    .C1(_07821_),
    .Y(_07824_));
 sky130_fd_sc_hd__a31oi_4 _18282_ (.A1(_07821_),
    .A2(net241),
    .A3(_07820_),
    .B1(_07810_),
    .Y(_07825_));
 sky130_fd_sc_hd__or4_2 _18283_ (.A(net259),
    .B(net256),
    .C(_07810_),
    .D(_07823_),
    .X(_07826_));
 sky130_fd_sc_hd__a311oi_4 _18284_ (.A1(_07821_),
    .A2(net241),
    .A3(_07820_),
    .B1(_07810_),
    .C1(_07899_),
    .Y(_07827_));
 sky130_fd_sc_hd__a2bb2oi_2 _18285_ (.A1_N(_07800_),
    .A2_N(_07822_),
    .B1(_07812_),
    .B2(_07824_),
    .Y(_07828_));
 sky130_fd_sc_hd__o21ai_1 _18286_ (.A1(_07810_),
    .A2(_07823_),
    .B1(_07899_),
    .Y(_07829_));
 sky130_fd_sc_hd__o32a_1 _18287_ (.A1(_06945_),
    .A2(_06967_),
    .A3(_07490_),
    .B1(_07497_),
    .B2(_07493_),
    .X(_07830_));
 sky130_fd_sc_hd__o32ai_4 _18288_ (.A1(_06945_),
    .A2(_06967_),
    .A3(_07490_),
    .B1(_07497_),
    .B2(_07493_),
    .Y(_07831_));
 sky130_fd_sc_hd__o21ai_1 _18289_ (.A1(_07888_),
    .A2(_07825_),
    .B1(_07830_),
    .Y(_07832_));
 sky130_fd_sc_hd__o21ai_1 _18290_ (.A1(_07827_),
    .A2(_07828_),
    .B1(_07831_),
    .Y(_07834_));
 sky130_fd_sc_hd__o21ai_1 _18291_ (.A1(_07827_),
    .A2(_07828_),
    .B1(_07830_),
    .Y(_07835_));
 sky130_fd_sc_hd__nand3b_1 _18292_ (.A_N(_07827_),
    .B(_07829_),
    .C(_07831_),
    .Y(_07836_));
 sky130_fd_sc_hd__o211ai_4 _18293_ (.A1(net259),
    .A2(net256),
    .B1(_07835_),
    .C1(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__or3_1 _18294_ (.A(net259),
    .B(net256),
    .C(_07825_),
    .X(_07838_));
 sky130_fd_sc_hd__o221ai_4 _18295_ (.A1(net259),
    .A2(net256),
    .B1(_07827_),
    .B2(_07832_),
    .C1(_07834_),
    .Y(_07839_));
 sky130_fd_sc_hd__o31a_2 _18296_ (.A1(_05996_),
    .A2(_07810_),
    .A3(_07823_),
    .B1(_07837_),
    .X(_07840_));
 sky130_fd_sc_hd__a21oi_2 _18297_ (.A1(_07507_),
    .A2(_07506_),
    .B1(_07503_),
    .Y(_07841_));
 sky130_fd_sc_hd__a21o_1 _18298_ (.A1(_07507_),
    .A2(_07506_),
    .B1(_07503_),
    .X(_07842_));
 sky130_fd_sc_hd__o221a_1 _18299_ (.A1(_06989_),
    .A2(net375),
    .B1(_05996_),
    .B2(_07825_),
    .C1(_07839_),
    .X(_07843_));
 sky130_fd_sc_hd__o221ai_4 _18300_ (.A1(_06989_),
    .A2(net375),
    .B1(_05996_),
    .B2(_07825_),
    .C1(_07839_),
    .Y(_07845_));
 sky130_fd_sc_hd__a2bb2oi_1 _18301_ (.A1_N(_06945_),
    .A2_N(_06967_),
    .B1(_07838_),
    .B2(_07839_),
    .Y(_07846_));
 sky130_fd_sc_hd__o211ai_4 _18302_ (.A1(_06945_),
    .A2(_06967_),
    .B1(_07826_),
    .C1(_07837_),
    .Y(_07847_));
 sky130_fd_sc_hd__a21oi_2 _18303_ (.A1(_07845_),
    .A2(_07847_),
    .B1(_07841_),
    .Y(_07848_));
 sky130_fd_sc_hd__a2bb2o_1 _18304_ (.A1_N(_07503_),
    .A2_N(_07509_),
    .B1(_07845_),
    .B2(_07847_),
    .X(_07849_));
 sky130_fd_sc_hd__a31oi_1 _18305_ (.A1(_07847_),
    .A2(_07841_),
    .A3(_07845_),
    .B1(_06294_),
    .Y(_07850_));
 sky130_fd_sc_hd__a31o_1 _18306_ (.A1(_07847_),
    .A2(_07841_),
    .A3(_07845_),
    .B1(_06294_),
    .X(_07851_));
 sky130_fd_sc_hd__a22o_1 _18307_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_07838_),
    .B2(_07839_),
    .X(_07852_));
 sky130_fd_sc_hd__a31o_1 _18308_ (.A1(_07044_),
    .A2(_07826_),
    .A3(_07837_),
    .B1(_07841_),
    .X(_07853_));
 sky130_fd_sc_hd__a21o_1 _18309_ (.A1(_07845_),
    .A2(_07847_),
    .B1(_07842_),
    .X(_07854_));
 sky130_fd_sc_hd__o221ai_2 _18310_ (.A1(_06291_),
    .A2(_06292_),
    .B1(_07843_),
    .B2(_07853_),
    .C1(_07854_),
    .Y(_07856_));
 sky130_fd_sc_hd__a2bb2oi_1 _18311_ (.A1_N(net212),
    .A2_N(_07840_),
    .B1(_07849_),
    .B2(_07850_),
    .Y(_07857_));
 sky130_fd_sc_hd__a2bb2o_1 _18312_ (.A1_N(net212),
    .A2_N(_07840_),
    .B1(_07849_),
    .B2(_07850_),
    .X(_07858_));
 sky130_fd_sc_hd__and3_1 _18313_ (.A(_06613_),
    .B(_07852_),
    .C(_07856_),
    .X(_07859_));
 sky130_fd_sc_hd__o221a_1 _18314_ (.A1(net212),
    .A2(_07840_),
    .B1(_07848_),
    .B2(_07851_),
    .C1(_06343_),
    .X(_07860_));
 sky130_fd_sc_hd__o221ai_4 _18315_ (.A1(net212),
    .A2(_07840_),
    .B1(_07848_),
    .B2(_07851_),
    .C1(_06343_),
    .Y(_07861_));
 sky130_fd_sc_hd__o211ai_2 _18316_ (.A1(net381),
    .A2(_06310_),
    .B1(_07852_),
    .C1(_07856_),
    .Y(_07862_));
 sky130_fd_sc_hd__o31a_1 _18317_ (.A1(_05862_),
    .A2(_07208_),
    .A3(_07514_),
    .B1(_07513_),
    .X(_07863_));
 sky130_fd_sc_hd__a221oi_2 _18318_ (.A1(_07206_),
    .A2(_07207_),
    .B1(_07513_),
    .B2(_05862_),
    .C1(_07208_),
    .Y(_07864_));
 sky130_fd_sc_hd__o2bb2ai_1 _18319_ (.A1_N(_07861_),
    .A2_N(_07862_),
    .B1(_07863_),
    .B2(_07518_),
    .Y(_07865_));
 sky130_fd_sc_hd__o211ai_2 _18320_ (.A1(_07525_),
    .A2(_07864_),
    .B1(_07862_),
    .C1(_07861_),
    .Y(_07867_));
 sky130_fd_sc_hd__o2bb2ai_1 _18321_ (.A1_N(_07861_),
    .A2_N(_07862_),
    .B1(_07864_),
    .B2(_07525_),
    .Y(_07868_));
 sky130_fd_sc_hd__o22ai_4 _18322_ (.A1(_07518_),
    .A2(_07863_),
    .B1(_06343_),
    .B2(_07857_),
    .Y(_07869_));
 sky130_fd_sc_hd__o221ai_2 _18323_ (.A1(_06608_),
    .A2(net237),
    .B1(_07860_),
    .B2(_07869_),
    .C1(_07868_),
    .Y(_07870_));
 sky130_fd_sc_hd__or3_1 _18324_ (.A(_06608_),
    .B(net237),
    .C(_07858_),
    .X(_07871_));
 sky130_fd_sc_hd__a31oi_2 _18325_ (.A1(_07865_),
    .A2(_07867_),
    .A3(_06612_),
    .B1(_07859_),
    .Y(_07872_));
 sky130_fd_sc_hd__a31o_1 _18326_ (.A1(_07865_),
    .A2(_07867_),
    .A3(_06612_),
    .B1(_07859_),
    .X(_07873_));
 sky130_fd_sc_hd__nand4_4 _18327_ (.A(_07218_),
    .B(_07222_),
    .C(_07522_),
    .D(_07524_),
    .Y(_07874_));
 sky130_fd_sc_hd__o211ai_4 _18328_ (.A1(_05545_),
    .A2(_07526_),
    .B1(_07532_),
    .C1(_07874_),
    .Y(_07875_));
 sky130_fd_sc_hd__and4_1 _18329_ (.A(_07529_),
    .B(_07532_),
    .C(_07874_),
    .D(_05851_),
    .X(_07876_));
 sky130_fd_sc_hd__o2111ai_2 _18330_ (.A1(_05545_),
    .A2(_07526_),
    .B1(_05851_),
    .C1(_07874_),
    .D1(_07532_),
    .Y(_07878_));
 sky130_fd_sc_hd__a31o_1 _18331_ (.A1(_07529_),
    .A2(_07532_),
    .A3(_07874_),
    .B1(_05851_),
    .X(_07879_));
 sky130_fd_sc_hd__a21oi_2 _18332_ (.A1(_05862_),
    .A2(_07875_),
    .B1(_06904_),
    .Y(_07880_));
 sky130_fd_sc_hd__o211ai_2 _18333_ (.A1(net230),
    .A2(_06901_),
    .B1(_07878_),
    .C1(_07879_),
    .Y(_07881_));
 sky130_fd_sc_hd__and3_1 _18334_ (.A(_07872_),
    .B(_07880_),
    .C(_07878_),
    .X(_07882_));
 sky130_fd_sc_hd__o211ai_4 _18335_ (.A1(_05862_),
    .A2(_07875_),
    .B1(_07880_),
    .C1(_07872_),
    .Y(_07883_));
 sky130_fd_sc_hd__o211a_1 _18336_ (.A1(_06612_),
    .A2(_07858_),
    .B1(_07870_),
    .C1(_07881_),
    .X(_07884_));
 sky130_fd_sc_hd__nand2_2 _18337_ (.A(_07873_),
    .B(_07881_),
    .Y(_07885_));
 sky130_fd_sc_hd__o32a_1 _18338_ (.A1(net407),
    .A2(_05218_),
    .A3(_07235_),
    .B1(_07534_),
    .B2(_07533_),
    .X(_07886_));
 sky130_fd_sc_hd__o32ai_4 _18339_ (.A1(net407),
    .A2(_05218_),
    .A3(_07235_),
    .B1(_07534_),
    .B2(_07533_),
    .Y(_07887_));
 sky130_fd_sc_hd__o211ai_2 _18340_ (.A1(_07533_),
    .A2(_07534_),
    .B1(_05545_),
    .C1(_07535_),
    .Y(_07889_));
 sky130_fd_sc_hd__o21ai_1 _18341_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_07887_),
    .Y(_07890_));
 sky130_fd_sc_hd__a22oi_4 _18342_ (.A1(_07228_),
    .A2(_07230_),
    .B1(_07887_),
    .B2(_05556_),
    .Y(_07891_));
 sky130_fd_sc_hd__a22oi_1 _18343_ (.A1(_07883_),
    .A2(_07885_),
    .B1(_07891_),
    .B2(_07889_),
    .Y(_07892_));
 sky130_fd_sc_hd__o2bb2ai_2 _18344_ (.A1_N(_07889_),
    .A2_N(_07891_),
    .B1(_07882_),
    .B2(_07884_),
    .Y(_07893_));
 sky130_fd_sc_hd__o2111a_1 _18345_ (.A1(_05556_),
    .A2(_07887_),
    .B1(_07885_),
    .C1(_07883_),
    .D1(_07891_),
    .X(_07894_));
 sky130_fd_sc_hd__o2111ai_4 _18346_ (.A1(_05556_),
    .A2(_07887_),
    .B1(_07885_),
    .C1(_07883_),
    .D1(_07891_),
    .Y(_07895_));
 sky130_fd_sc_hd__nand2_1 _18347_ (.A(_07893_),
    .B(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__nand3_4 _18348_ (.A(_07893_),
    .B(_07895_),
    .C(_05239_),
    .Y(_07897_));
 sky130_fd_sc_hd__inv_2 _18349_ (.A(_07897_),
    .Y(_07898_));
 sky130_fd_sc_hd__a21oi_2 _18350_ (.A1(_07893_),
    .A2(_07895_),
    .B1(_05239_),
    .Y(_07900_));
 sky130_fd_sc_hd__o21ai_1 _18351_ (.A1(_07892_),
    .A2(_07894_),
    .B1(_05250_),
    .Y(_07901_));
 sky130_fd_sc_hd__a2bb2o_1 _18352_ (.A1_N(_03289_),
    .A2_N(_07539_),
    .B1(_07897_),
    .B2(_07901_),
    .X(_07902_));
 sky130_fd_sc_hd__a21oi_1 _18353_ (.A1(_05250_),
    .A2(_07896_),
    .B1(_07541_),
    .Y(_07903_));
 sky130_fd_sc_hd__nand2_1 _18354_ (.A(_07901_),
    .B(_07540_),
    .Y(_07904_));
 sky130_fd_sc_hd__a31oi_1 _18355_ (.A1(_07901_),
    .A2(_07540_),
    .A3(_07897_),
    .B1(_07550_),
    .Y(_07905_));
 sky130_fd_sc_hd__a2bb2o_1 _18356_ (.A1_N(net163),
    .A2_N(_07896_),
    .B1(_07902_),
    .B2(_07905_),
    .X(_07906_));
 sky130_fd_sc_hd__o2bb2a_1 _18357_ (.A1_N(_07905_),
    .A2_N(_07902_),
    .B1(_07896_),
    .B2(net163),
    .X(_07907_));
 sky130_fd_sc_hd__o31ai_4 _18358_ (.A1(net45),
    .A2(net46),
    .A3(_07226_),
    .B1(net409),
    .Y(_07908_));
 sky130_fd_sc_hd__o311a_4 _18359_ (.A1(net45),
    .A2(net46),
    .A3(_07226_),
    .B1(net47),
    .C1(net409),
    .X(_07909_));
 sky130_fd_sc_hd__and2b_4 _18360_ (.A_N(net47),
    .B(_07908_),
    .X(_07911_));
 sky130_fd_sc_hd__nor2_8 _18361_ (.A(net47),
    .B(_07908_),
    .Y(_07912_));
 sky130_fd_sc_hd__clkinv_4 _18362_ (.A(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__and2_4 _18363_ (.A(_07908_),
    .B(net47),
    .X(_07914_));
 sky130_fd_sc_hd__clkinv_4 _18364_ (.A(_07914_),
    .Y(_07915_));
 sky130_fd_sc_hd__nor2_8 _18365_ (.A(_07909_),
    .B(_07911_),
    .Y(_07916_));
 sky130_fd_sc_hd__nor2_8 _18366_ (.A(_07912_),
    .B(_07914_),
    .Y(_07917_));
 sky130_fd_sc_hd__o21ai_1 _18367_ (.A1(_03289_),
    .A2(_07917_),
    .B1(_07907_),
    .Y(_07918_));
 sky130_fd_sc_hd__nand2_1 _18368_ (.A(net1),
    .B(_07906_),
    .Y(_07919_));
 sky130_fd_sc_hd__o31a_1 _18369_ (.A1(_03289_),
    .A2(_07907_),
    .A3(_07917_),
    .B1(_07918_),
    .X(_07920_));
 sky130_fd_sc_hd__and3_1 _18370_ (.A(_07920_),
    .B(_07553_),
    .C(_05119_),
    .X(_07922_));
 sky130_fd_sc_hd__a21oi_1 _18371_ (.A1(_05119_),
    .A2(_07553_),
    .B1(_07920_),
    .Y(_07923_));
 sky130_fd_sc_hd__nor2_1 _18372_ (.A(_07922_),
    .B(_07923_),
    .Y(net79));
 sky130_fd_sc_hd__o22a_1 _18373_ (.A1(_04832_),
    .A2(_04942_),
    .B1(_07553_),
    .B2(_07920_),
    .X(_07924_));
 sky130_fd_sc_hd__o21ai_2 _18374_ (.A1(_06332_),
    .A2(_07858_),
    .B1(_07869_),
    .Y(_07925_));
 sky130_fd_sc_hd__or4_4 _18375_ (.A(net13),
    .B(net14),
    .C(net15),
    .D(_06913_),
    .X(_07926_));
 sky130_fd_sc_hd__o21ai_4 _18376_ (.A1(net15),
    .A2(_07554_),
    .B1(net410),
    .Y(_07927_));
 sky130_fd_sc_hd__nor2_8 _18377_ (.A(net16),
    .B(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__or3b_4 _18378_ (.A(_03399_),
    .B(net16),
    .C_N(_07926_),
    .X(_07929_));
 sky130_fd_sc_hd__and2_4 _18379_ (.A(_07927_),
    .B(net16),
    .X(_07930_));
 sky130_fd_sc_hd__nand2_8 _18380_ (.A(_07927_),
    .B(net16),
    .Y(_07932_));
 sky130_fd_sc_hd__o211ai_4 _18381_ (.A1(net15),
    .A2(_07554_),
    .B1(net16),
    .C1(net410),
    .Y(_07933_));
 sky130_fd_sc_hd__a21o_4 _18382_ (.A1(_07926_),
    .A2(net410),
    .B1(net16),
    .X(_07934_));
 sky130_fd_sc_hd__nand2_8 _18383_ (.A(_07933_),
    .B(_07934_),
    .Y(_07935_));
 sky130_fd_sc_hd__nand2_8 _18384_ (.A(_07929_),
    .B(_07932_),
    .Y(_07936_));
 sky130_fd_sc_hd__and3_1 _18385_ (.A(_07934_),
    .B(net33),
    .C(_07933_),
    .X(_07937_));
 sky130_fd_sc_hd__o21ai_1 _18386_ (.A1(_07928_),
    .A2(_07930_),
    .B1(net33),
    .Y(_07938_));
 sky130_fd_sc_hd__o22a_2 _18387_ (.A1(_05130_),
    .A2(_05152_),
    .B1(_03178_),
    .B2(_07935_),
    .X(_07939_));
 sky130_fd_sc_hd__a31o_2 _18388_ (.A1(_07934_),
    .A2(net33),
    .A3(_07933_),
    .B1(net405),
    .X(_07940_));
 sky130_fd_sc_hd__a31o_1 _18389_ (.A1(net33),
    .A2(_07933_),
    .A3(_07934_),
    .B1(net202),
    .X(_07941_));
 sky130_fd_sc_hd__o21ai_2 _18390_ (.A1(_07566_),
    .A2(_07935_),
    .B1(_07941_),
    .Y(_07943_));
 sky130_fd_sc_hd__a21o_1 _18391_ (.A1(_07569_),
    .A2(_07573_),
    .B1(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__o211ai_2 _18392_ (.A1(_07564_),
    .A2(_07249_),
    .B1(_07943_),
    .C1(_07573_),
    .Y(_07945_));
 sky130_fd_sc_hd__a21oi_2 _18393_ (.A1(_07944_),
    .A2(_07945_),
    .B1(_05185_),
    .Y(_07946_));
 sky130_fd_sc_hd__a21o_1 _18394_ (.A1(_07944_),
    .A2(_07945_),
    .B1(_05185_),
    .X(_07947_));
 sky130_fd_sc_hd__or4_1 _18395_ (.A(_05348_),
    .B(net401),
    .C(_07939_),
    .D(_07946_),
    .X(_07948_));
 sky130_fd_sc_hd__o21ai_1 _18396_ (.A1(_07939_),
    .A2(_07946_),
    .B1(net224),
    .Y(_07949_));
 sky130_fd_sc_hd__o21a_1 _18397_ (.A1(_07242_),
    .A2(_07243_),
    .B1(_07947_),
    .X(_07950_));
 sky130_fd_sc_hd__or3_1 _18398_ (.A(_07244_),
    .B(_07245_),
    .C(_07946_),
    .X(_07951_));
 sky130_fd_sc_hd__o221ai_1 _18399_ (.A1(_07242_),
    .A2(_07243_),
    .B1(_07937_),
    .B2(net405),
    .C1(_07947_),
    .Y(_07952_));
 sky130_fd_sc_hd__o41a_4 _18400_ (.A1(_07244_),
    .A2(_07245_),
    .A3(_07939_),
    .A4(_07946_),
    .B1(_07949_),
    .X(_07954_));
 sky130_fd_sc_hd__o22ai_2 _18401_ (.A1(net227),
    .A2(_07577_),
    .B1(_07588_),
    .B2(_07591_),
    .Y(_07955_));
 sky130_fd_sc_hd__o21ai_1 _18402_ (.A1(_07586_),
    .A2(_07587_),
    .B1(_07583_),
    .Y(_07956_));
 sky130_fd_sc_hd__o21bai_2 _18403_ (.A1(_07956_),
    .A2(_07591_),
    .B1_N(_07579_),
    .Y(_07957_));
 sky130_fd_sc_hd__o211ai_4 _18404_ (.A1(net225),
    .A2(_07576_),
    .B1(_07954_),
    .C1(_07955_),
    .Y(_07958_));
 sky130_fd_sc_hd__a21oi_1 _18405_ (.A1(_07949_),
    .A2(_07952_),
    .B1(_07579_),
    .Y(_07959_));
 sky130_fd_sc_hd__nand2_1 _18406_ (.A(_07597_),
    .B(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__a21oi_1 _18407_ (.A1(_07597_),
    .A2(_07959_),
    .B1(_05392_),
    .Y(_07961_));
 sky130_fd_sc_hd__o211ai_2 _18408_ (.A1(_05348_),
    .A2(net401),
    .B1(_07958_),
    .C1(_07960_),
    .Y(_07962_));
 sky130_fd_sc_hd__a32oi_4 _18409_ (.A1(_05392_),
    .A2(_07940_),
    .A3(_07947_),
    .B1(_07961_),
    .B2(_07958_),
    .Y(_07963_));
 sky130_fd_sc_hd__or3_2 _18410_ (.A(_05676_),
    .B(_05698_),
    .C(_07963_),
    .X(_07965_));
 sky130_fd_sc_hd__inv_2 _18411_ (.A(_07965_),
    .Y(_07966_));
 sky130_fd_sc_hd__a2bb2oi_1 _18412_ (.A1_N(_06914_),
    .A2_N(_06916_),
    .B1(_07948_),
    .B2(_07962_),
    .Y(_07967_));
 sky130_fd_sc_hd__a22o_1 _18413_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_07948_),
    .B2(_07962_),
    .X(_07968_));
 sky130_fd_sc_hd__o311a_1 _18414_ (.A1(_05403_),
    .A2(_07939_),
    .A3(_07946_),
    .B1(net227),
    .C1(_07962_),
    .X(_07969_));
 sky130_fd_sc_hd__o21ai_1 _18415_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_07963_),
    .Y(_07970_));
 sky130_fd_sc_hd__nor2_2 _18416_ (.A(_07967_),
    .B(_07969_),
    .Y(_07971_));
 sky130_fd_sc_hd__o211ai_2 _18417_ (.A1(_06950_),
    .A2(_06958_),
    .B1(_06662_),
    .C1(_06955_),
    .Y(_07972_));
 sky130_fd_sc_hd__a211oi_2 _18418_ (.A1(_07261_),
    .A2(_07278_),
    .B1(_07972_),
    .C1(_07277_),
    .Y(_07973_));
 sky130_fd_sc_hd__o21ai_1 _18419_ (.A1(net232),
    .A2(_07600_),
    .B1(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__a21oi_1 _18420_ (.A1(_07973_),
    .A2(_07606_),
    .B1(_07601_),
    .Y(_07976_));
 sky130_fd_sc_hd__o211a_2 _18421_ (.A1(_07605_),
    .A2(_07609_),
    .B1(_07974_),
    .C1(_07602_),
    .X(_07977_));
 sky130_fd_sc_hd__o211ai_2 _18422_ (.A1(_07605_),
    .A2(_07609_),
    .B1(_07974_),
    .C1(_07602_),
    .Y(_07978_));
 sky130_fd_sc_hd__nor4_1 _18423_ (.A(_06671_),
    .B(_07277_),
    .C(_07972_),
    .D(_07279_),
    .Y(_07979_));
 sky130_fd_sc_hd__nand4_2 _18424_ (.A(_07602_),
    .B(_07973_),
    .C(_07606_),
    .D(_06673_),
    .Y(_07980_));
 sky130_fd_sc_hd__a22oi_4 _18425_ (.A1(_07607_),
    .A2(_07979_),
    .B1(_07610_),
    .B2(_07976_),
    .Y(_07981_));
 sky130_fd_sc_hd__a31o_1 _18426_ (.A1(_06673_),
    .A2(_07607_),
    .A3(_07973_),
    .B1(_07977_),
    .X(_07982_));
 sky130_fd_sc_hd__nand3_2 _18427_ (.A(_07968_),
    .B(_07970_),
    .C(_07980_),
    .Y(_07983_));
 sky130_fd_sc_hd__o311a_1 _18428_ (.A1(_06671_),
    .A2(_07601_),
    .A3(_07974_),
    .B1(_07978_),
    .C1(_07971_),
    .X(_07984_));
 sky130_fd_sc_hd__nand3_2 _18429_ (.A(_07971_),
    .B(_07978_),
    .C(_07980_),
    .Y(_07985_));
 sky130_fd_sc_hd__o22ai_1 _18430_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_07971_),
    .B2(_07981_),
    .Y(_07987_));
 sky130_fd_sc_hd__o221a_1 _18431_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_07971_),
    .B2(_07981_),
    .C1(_07985_),
    .X(_07988_));
 sky130_fd_sc_hd__o221ai_4 _18432_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_07971_),
    .B2(_07981_),
    .C1(_07985_),
    .Y(_07989_));
 sky130_fd_sc_hd__o22a_1 _18433_ (.A1(net359),
    .A2(_07963_),
    .B1(_07984_),
    .B2(_07987_),
    .X(_07990_));
 sky130_fd_sc_hd__o211a_2 _18434_ (.A1(_07966_),
    .A2(_07988_),
    .B1(_06804_),
    .C1(_06826_),
    .X(_07991_));
 sky130_fd_sc_hd__or3_4 _18435_ (.A(_06793_),
    .B(_06815_),
    .C(_07990_),
    .X(_07992_));
 sky130_fd_sc_hd__o221ai_4 _18436_ (.A1(net254),
    .A2(_07290_),
    .B1(_07299_),
    .B2(_07301_),
    .C1(_07618_),
    .Y(_07993_));
 sky130_fd_sc_hd__o22ai_4 _18437_ (.A1(_07613_),
    .A2(_07620_),
    .B1(_07617_),
    .B2(_07626_),
    .Y(_07994_));
 sky130_fd_sc_hd__o22a_1 _18438_ (.A1(_06626_),
    .A2(_06627_),
    .B1(_07984_),
    .B2(_07987_),
    .X(_07995_));
 sky130_fd_sc_hd__o211a_2 _18439_ (.A1(net359),
    .A2(_07963_),
    .B1(net234),
    .C1(_07989_),
    .X(_07996_));
 sky130_fd_sc_hd__o211ai_4 _18440_ (.A1(net359),
    .A2(_07963_),
    .B1(net234),
    .C1(_07989_),
    .Y(_07998_));
 sky130_fd_sc_hd__a2bb2oi_4 _18441_ (.A1_N(_06622_),
    .A2_N(_06624_),
    .B1(_07965_),
    .B2(_07989_),
    .Y(_07999_));
 sky130_fd_sc_hd__o22ai_4 _18442_ (.A1(_06622_),
    .A2(_06624_),
    .B1(_07966_),
    .B2(_07988_),
    .Y(_08000_));
 sky130_fd_sc_hd__a21oi_1 _18443_ (.A1(_07995_),
    .A2(_07965_),
    .B1(_07999_),
    .Y(_08001_));
 sky130_fd_sc_hd__nand4_4 _18444_ (.A(_07622_),
    .B(_07993_),
    .C(_07998_),
    .D(_08000_),
    .Y(_08002_));
 sky130_fd_sc_hd__o21ai_4 _18445_ (.A1(_07996_),
    .A2(_07999_),
    .B1(_07994_),
    .Y(_08003_));
 sky130_fd_sc_hd__o211a_1 _18446_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_08002_),
    .C1(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__o211ai_4 _18447_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_08002_),
    .C1(_08003_),
    .Y(_08005_));
 sky130_fd_sc_hd__a31o_2 _18448_ (.A1(_08003_),
    .A2(net357),
    .A3(_08002_),
    .B1(_07991_),
    .X(_08006_));
 sky130_fd_sc_hd__a2bb2oi_4 _18449_ (.A1_N(_06305_),
    .A2_N(net283),
    .B1(_07992_),
    .B2(_08005_),
    .Y(_08007_));
 sky130_fd_sc_hd__o22ai_4 _18450_ (.A1(_06305_),
    .A2(net283),
    .B1(_07991_),
    .B2(_08004_),
    .Y(_08009_));
 sky130_fd_sc_hd__a31oi_2 _18451_ (.A1(_08002_),
    .A2(_08003_),
    .A3(net357),
    .B1(net251),
    .Y(_08010_));
 sky130_fd_sc_hd__o211a_1 _18452_ (.A1(net357),
    .A2(_07990_),
    .B1(_06314_),
    .C1(_08005_),
    .X(_08011_));
 sky130_fd_sc_hd__o211ai_2 _18453_ (.A1(net357),
    .A2(_07990_),
    .B1(_06314_),
    .C1(_08005_),
    .Y(_08012_));
 sky130_fd_sc_hd__a21oi_1 _18454_ (.A1(_07992_),
    .A2(_08010_),
    .B1(_08007_),
    .Y(_08013_));
 sky130_fd_sc_hd__a21oi_2 _18455_ (.A1(_07640_),
    .A2(_07639_),
    .B1(_07635_),
    .Y(_08014_));
 sky130_fd_sc_hd__o21bai_2 _18456_ (.A1(_07638_),
    .A2(_07641_),
    .B1_N(_07635_),
    .Y(_08015_));
 sky130_fd_sc_hd__a21oi_1 _18457_ (.A1(_08009_),
    .A2(_08012_),
    .B1(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__o21ai_2 _18458_ (.A1(_08007_),
    .A2(_08011_),
    .B1(_08014_),
    .Y(_08017_));
 sky130_fd_sc_hd__a211oi_2 _18459_ (.A1(_08010_),
    .A2(_07992_),
    .B1(_08007_),
    .C1(_08014_),
    .Y(_08018_));
 sky130_fd_sc_hd__nand3_1 _18460_ (.A(_08009_),
    .B(_08012_),
    .C(_08015_),
    .Y(_08020_));
 sky130_fd_sc_hd__o22ai_4 _18461_ (.A1(net373),
    .A2(net371),
    .B1(_08016_),
    .B2(_08018_),
    .Y(_08021_));
 sky130_fd_sc_hd__a21oi_2 _18462_ (.A1(_07992_),
    .A2(_08005_),
    .B1(net355),
    .Y(_08022_));
 sky130_fd_sc_hd__a211o_1 _18463_ (.A1(_07992_),
    .A2(_08005_),
    .B1(net373),
    .C1(net371),
    .X(_08023_));
 sky130_fd_sc_hd__nand3_1 _18464_ (.A(_08017_),
    .B(_08020_),
    .C(net355),
    .Y(_08024_));
 sky130_fd_sc_hd__a31o_2 _18465_ (.A1(_08017_),
    .A2(_08020_),
    .A3(net355),
    .B1(_08022_),
    .X(_08025_));
 sky130_fd_sc_hd__a2bb2oi_1 _18466_ (.A1_N(_06009_),
    .A2_N(_06010_),
    .B1(_08023_),
    .B2(_08024_),
    .Y(_08026_));
 sky130_fd_sc_hd__o211ai_4 _18467_ (.A1(_08006_),
    .A2(net355),
    .B1(net253),
    .C1(_08021_),
    .Y(_08027_));
 sky130_fd_sc_hd__a31o_1 _18468_ (.A1(_08017_),
    .A2(_08020_),
    .A3(net355),
    .B1(net253),
    .X(_08028_));
 sky130_fd_sc_hd__and3_1 _18469_ (.A(_08024_),
    .B(net254),
    .C(_08023_),
    .X(_08029_));
 sky130_fd_sc_hd__a311o_2 _18470_ (.A1(_08017_),
    .A2(_08020_),
    .A3(net355),
    .B1(_08022_),
    .C1(net253),
    .X(_08031_));
 sky130_fd_sc_hd__o2bb2ai_2 _18471_ (.A1_N(net262),
    .A2_N(_07649_),
    .B1(_07657_),
    .B2(_07328_),
    .Y(_08032_));
 sky130_fd_sc_hd__o22ai_2 _18472_ (.A1(net262),
    .A2(_07649_),
    .B1(_08032_),
    .B2(_07662_),
    .Y(_08033_));
 sky130_fd_sc_hd__nand4_2 _18473_ (.A(_07654_),
    .B(_07665_),
    .C(_08027_),
    .D(_08031_),
    .Y(_08034_));
 sky130_fd_sc_hd__o21ai_1 _18474_ (.A1(_08026_),
    .A2(_08029_),
    .B1(_08033_),
    .Y(_08035_));
 sky130_fd_sc_hd__o211ai_4 _18475_ (.A1(net353),
    .A2(net352),
    .B1(_08034_),
    .C1(_08035_),
    .Y(_08036_));
 sky130_fd_sc_hd__o311a_1 _18476_ (.A1(_07691_),
    .A2(_08006_),
    .A3(net371),
    .B1(_08732_),
    .C1(_08021_),
    .X(_08037_));
 sky130_fd_sc_hd__o211ai_2 _18477_ (.A1(_08026_),
    .A2(_08029_),
    .B1(_07654_),
    .C1(_07665_),
    .Y(_08038_));
 sky130_fd_sc_hd__nand3_1 _18478_ (.A(_08033_),
    .B(_08031_),
    .C(_08027_),
    .Y(_08039_));
 sky130_fd_sc_hd__o211ai_1 _18479_ (.A1(net353),
    .A2(_08700_),
    .B1(_08038_),
    .C1(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__o21ai_4 _18480_ (.A1(net338),
    .A2(_08025_),
    .B1(_08036_),
    .Y(_08042_));
 sky130_fd_sc_hd__inv_2 _18481_ (.A(_08042_),
    .Y(_08043_));
 sky130_fd_sc_hd__o211a_1 _18482_ (.A1(net338),
    .A2(_08025_),
    .B1(_08036_),
    .C1(net261),
    .X(_08044_));
 sky130_fd_sc_hd__o211ai_4 _18483_ (.A1(net338),
    .A2(_08025_),
    .B1(_08036_),
    .C1(net261),
    .Y(_08045_));
 sky130_fd_sc_hd__a31o_1 _18484_ (.A1(_08038_),
    .A2(_08039_),
    .A3(net338),
    .B1(net261),
    .X(_08046_));
 sky130_fd_sc_hd__nand3b_2 _18485_ (.A_N(_08037_),
    .B(_08040_),
    .C(net262),
    .Y(_08047_));
 sky130_fd_sc_hd__o21a_1 _18486_ (.A1(_08037_),
    .A2(_08046_),
    .B1(_08045_),
    .X(_08048_));
 sky130_fd_sc_hd__nand3_1 _18487_ (.A(_07041_),
    .B(_07043_),
    .C(_06730_),
    .Y(_08049_));
 sky130_fd_sc_hd__nor3_2 _18488_ (.A(_07343_),
    .B(_08049_),
    .C(_07345_),
    .Y(_08050_));
 sky130_fd_sc_hd__nand2_1 _18489_ (.A(_08050_),
    .B(_07677_),
    .Y(_08051_));
 sky130_fd_sc_hd__a21oi_1 _18490_ (.A1(_08050_),
    .A2(_07677_),
    .B1(_07678_),
    .Y(_08053_));
 sky130_fd_sc_hd__o211ai_4 _18491_ (.A1(_07683_),
    .A2(_07676_),
    .B1(_07679_),
    .C1(_08051_),
    .Y(_08054_));
 sky130_fd_sc_hd__o211ai_1 _18492_ (.A1(_06443_),
    .A2(_06723_),
    .B1(_08050_),
    .C1(_07679_),
    .Y(_08055_));
 sky130_fd_sc_hd__nand4b_4 _18493_ (.A_N(_06724_),
    .B(_07677_),
    .C(_07679_),
    .D(_08050_),
    .Y(_08056_));
 sky130_fd_sc_hd__a2bb2oi_1 _18494_ (.A1_N(_07676_),
    .A2_N(_08055_),
    .B1(_07685_),
    .B2(_08053_),
    .Y(_08057_));
 sky130_fd_sc_hd__o211ai_1 _18495_ (.A1(_08037_),
    .A2(_08046_),
    .B1(_08056_),
    .C1(_08045_),
    .Y(_08058_));
 sky130_fd_sc_hd__a21oi_1 _18496_ (.A1(_07685_),
    .A2(_08053_),
    .B1(_08058_),
    .Y(_08059_));
 sky130_fd_sc_hd__nand4_4 _18497_ (.A(_08045_),
    .B(_08047_),
    .C(_08054_),
    .D(_08056_),
    .Y(_08060_));
 sky130_fd_sc_hd__a22o_2 _18498_ (.A1(_08045_),
    .A2(_08047_),
    .B1(_08054_),
    .B2(_08056_),
    .X(_08061_));
 sky130_fd_sc_hd__o22ai_1 _18499_ (.A1(_09785_),
    .A2(net349),
    .B1(_08048_),
    .B2(_08057_),
    .Y(_08062_));
 sky130_fd_sc_hd__nand3_2 _18500_ (.A(_08061_),
    .B(net336),
    .C(_08060_),
    .Y(_08064_));
 sky130_fd_sc_hd__o211a_2 _18501_ (.A1(net338),
    .A2(_08025_),
    .B1(_08036_),
    .C1(_09840_),
    .X(_08065_));
 sky130_fd_sc_hd__or3_2 _18502_ (.A(_09785_),
    .B(net349),
    .C(_08042_),
    .X(_08066_));
 sky130_fd_sc_hd__a31oi_4 _18503_ (.A1(_08061_),
    .A2(net336),
    .A3(_08060_),
    .B1(_08065_),
    .Y(_08067_));
 sky130_fd_sc_hd__o22ai_2 _18504_ (.A1(net336),
    .A2(_08042_),
    .B1(_08059_),
    .B2(_08062_),
    .Y(_08068_));
 sky130_fd_sc_hd__a21oi_2 _18505_ (.A1(_08064_),
    .A2(_08066_),
    .B1(net333),
    .Y(_08069_));
 sky130_fd_sc_hd__or3_2 _18506_ (.A(_11046_),
    .B(_11057_),
    .C(_08067_),
    .X(_08070_));
 sky130_fd_sc_hd__a31o_1 _18507_ (.A1(_08061_),
    .A2(net336),
    .A3(_08060_),
    .B1(net291),
    .X(_08071_));
 sky130_fd_sc_hd__a311oi_4 _18508_ (.A1(_08061_),
    .A2(net336),
    .A3(_08060_),
    .B1(_08065_),
    .C1(net291),
    .Y(_08072_));
 sky130_fd_sc_hd__nand3_2 _18509_ (.A(_08064_),
    .B(_08066_),
    .C(net267),
    .Y(_08073_));
 sky130_fd_sc_hd__a22oi_4 _18510_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_08064_),
    .B2(_08066_),
    .Y(_08075_));
 sky130_fd_sc_hd__o21ai_4 _18511_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_08068_),
    .Y(_08076_));
 sky130_fd_sc_hd__a21o_1 _18512_ (.A1(_07693_),
    .A2(_07696_),
    .B1(_07697_),
    .X(_08077_));
 sky130_fd_sc_hd__a21oi_2 _18513_ (.A1(_07693_),
    .A2(_07696_),
    .B1(_07697_),
    .Y(_08078_));
 sky130_fd_sc_hd__o21a_1 _18514_ (.A1(_08072_),
    .A2(_08075_),
    .B1(_08078_),
    .X(_08079_));
 sky130_fd_sc_hd__o21bai_4 _18515_ (.A1(_08072_),
    .A2(_08075_),
    .B1_N(_08077_),
    .Y(_08080_));
 sky130_fd_sc_hd__o21ai_2 _18516_ (.A1(net267),
    .A2(_08067_),
    .B1(_08077_),
    .Y(_08081_));
 sky130_fd_sc_hd__o211ai_4 _18517_ (.A1(_08065_),
    .A2(_08071_),
    .B1(_08077_),
    .C1(_08076_),
    .Y(_08082_));
 sky130_fd_sc_hd__o22ai_2 _18518_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_08072_),
    .B2(_08081_),
    .Y(_08083_));
 sky130_fd_sc_hd__o211ai_4 _18519_ (.A1(_08072_),
    .A2(_08081_),
    .B1(net333),
    .C1(_08080_),
    .Y(_08084_));
 sky130_fd_sc_hd__a31oi_4 _18520_ (.A1(_08080_),
    .A2(_08082_),
    .A3(net333),
    .B1(_08069_),
    .Y(_08086_));
 sky130_fd_sc_hd__o22ai_4 _18521_ (.A1(net333),
    .A2(_08067_),
    .B1(_08079_),
    .B2(_08083_),
    .Y(_08087_));
 sky130_fd_sc_hd__o2bb2a_1 _18522_ (.A1_N(net298),
    .A2_N(_07707_),
    .B1(_07712_),
    .B2(_07381_),
    .X(_08088_));
 sky130_fd_sc_hd__o221a_1 _18523_ (.A1(_07377_),
    .A2(_07379_),
    .B1(net298),
    .B2(_07707_),
    .C1(_07382_),
    .X(_08089_));
 sky130_fd_sc_hd__o32a_1 _18524_ (.A1(net339),
    .A2(_04184_),
    .A3(_07707_),
    .B1(_07710_),
    .B2(_07714_),
    .X(_08090_));
 sky130_fd_sc_hd__a31oi_1 _18525_ (.A1(_08080_),
    .A2(_08082_),
    .A3(net333),
    .B1(net293),
    .Y(_08091_));
 sky130_fd_sc_hd__a311oi_4 _18526_ (.A1(_08080_),
    .A2(_08082_),
    .A3(net333),
    .B1(net293),
    .C1(_08069_),
    .Y(_08092_));
 sky130_fd_sc_hd__o211ai_4 _18527_ (.A1(net333),
    .A2(_08067_),
    .B1(net295),
    .C1(_08084_),
    .Y(_08093_));
 sky130_fd_sc_hd__a2bb2oi_4 _18528_ (.A1_N(_05242_),
    .A2_N(net314),
    .B1(_08070_),
    .B2(_08084_),
    .Y(_08094_));
 sky130_fd_sc_hd__a22o_1 _18529_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_08070_),
    .B2(_08084_),
    .X(_08095_));
 sky130_fd_sc_hd__o211ai_1 _18530_ (.A1(_07708_),
    .A2(_08088_),
    .B1(_08093_),
    .C1(_08095_),
    .Y(_08097_));
 sky130_fd_sc_hd__o22ai_1 _18531_ (.A1(_07710_),
    .A2(_08089_),
    .B1(_08092_),
    .B2(_08094_),
    .Y(_08098_));
 sky130_fd_sc_hd__o21ai_1 _18532_ (.A1(net295),
    .A2(_08086_),
    .B1(_08090_),
    .Y(_08099_));
 sky130_fd_sc_hd__o211ai_4 _18533_ (.A1(_07710_),
    .A2(_08089_),
    .B1(_08093_),
    .C1(_08095_),
    .Y(_08100_));
 sky130_fd_sc_hd__o22ai_4 _18534_ (.A1(_07708_),
    .A2(_08088_),
    .B1(_08092_),
    .B2(_08094_),
    .Y(_08101_));
 sky130_fd_sc_hd__nand3_2 _18535_ (.A(_08097_),
    .B(_08098_),
    .C(net312),
    .Y(_08102_));
 sky130_fd_sc_hd__a21oi_1 _18536_ (.A1(_08070_),
    .A2(_08084_),
    .B1(net312),
    .Y(_08103_));
 sky130_fd_sc_hd__or3_1 _18537_ (.A(_12670_),
    .B(_12681_),
    .C(_08086_),
    .X(_08104_));
 sky130_fd_sc_hd__o221ai_4 _18538_ (.A1(_12670_),
    .A2(_12681_),
    .B1(_08092_),
    .B2(_08099_),
    .C1(_08101_),
    .Y(_08105_));
 sky130_fd_sc_hd__a31oi_4 _18539_ (.A1(_08100_),
    .A2(_08101_),
    .A3(net312),
    .B1(_08103_),
    .Y(_08106_));
 sky130_fd_sc_hd__a31oi_2 _18540_ (.A1(_08100_),
    .A2(_08101_),
    .A3(net312),
    .B1(net298),
    .Y(_08108_));
 sky130_fd_sc_hd__and3_1 _18541_ (.A(_08105_),
    .B(net299),
    .C(_08104_),
    .X(_08109_));
 sky130_fd_sc_hd__o211ai_4 _18542_ (.A1(net312),
    .A2(_08086_),
    .B1(net299),
    .C1(_08105_),
    .Y(_08110_));
 sky130_fd_sc_hd__a22oi_1 _18543_ (.A1(_04173_),
    .A2(_04195_),
    .B1(_08104_),
    .B2(_08105_),
    .Y(_08111_));
 sky130_fd_sc_hd__o211ai_4 _18544_ (.A1(_08087_),
    .A2(net312),
    .B1(net298),
    .C1(_08102_),
    .Y(_08112_));
 sky130_fd_sc_hd__a21oi_1 _18545_ (.A1(_07732_),
    .A2(_07734_),
    .B1(_07721_),
    .Y(_08113_));
 sky130_fd_sc_hd__a31oi_2 _18546_ (.A1(_07725_),
    .A2(_07732_),
    .A3(_07734_),
    .B1(_07721_),
    .Y(_08114_));
 sky130_fd_sc_hd__o22ai_2 _18547_ (.A1(_02137_),
    .A2(_07720_),
    .B1(_07737_),
    .B2(_07731_),
    .Y(_08115_));
 sky130_fd_sc_hd__o2bb2ai_2 _18548_ (.A1_N(_08110_),
    .A2_N(_08112_),
    .B1(_08113_),
    .B2(_07723_),
    .Y(_08116_));
 sky130_fd_sc_hd__nand3_2 _18549_ (.A(_08110_),
    .B(_08112_),
    .C(_08115_),
    .Y(_08117_));
 sky130_fd_sc_hd__o211a_1 _18550_ (.A1(_08087_),
    .A2(net312),
    .B1(_00066_),
    .C1(_08102_),
    .X(_08119_));
 sky130_fd_sc_hd__or3_1 _18551_ (.A(net324),
    .B(_00033_),
    .C(_08106_),
    .X(_08120_));
 sky130_fd_sc_hd__nand3_1 _18552_ (.A(_08116_),
    .B(_08117_),
    .C(net309),
    .Y(_08121_));
 sky130_fd_sc_hd__a31o_1 _18553_ (.A1(_08116_),
    .A2(_08117_),
    .A3(net309),
    .B1(_08119_),
    .X(_08122_));
 sky130_fd_sc_hd__a2bb2oi_1 _18554_ (.A1_N(_02049_),
    .A2_N(net342),
    .B1(_08120_),
    .B2(_08121_),
    .Y(_08123_));
 sky130_fd_sc_hd__o21ai_2 _18555_ (.A1(_02049_),
    .A2(net342),
    .B1(_08122_),
    .Y(_08124_));
 sky130_fd_sc_hd__o211a_1 _18556_ (.A1(net309),
    .A2(_08106_),
    .B1(_02137_),
    .C1(_08121_),
    .X(_08125_));
 sky130_fd_sc_hd__a311o_1 _18557_ (.A1(_08116_),
    .A2(_08117_),
    .A3(net309),
    .B1(_08119_),
    .C1(_02148_),
    .X(_08126_));
 sky130_fd_sc_hd__o22a_1 _18558_ (.A1(_07748_),
    .A2(_07742_),
    .B1(_07752_),
    .B2(_07750_),
    .X(_08127_));
 sky130_fd_sc_hd__o22ai_4 _18559_ (.A1(_07748_),
    .A2(_07742_),
    .B1(_07752_),
    .B2(_07750_),
    .Y(_08128_));
 sky130_fd_sc_hd__o21a_1 _18560_ (.A1(_02148_),
    .A2(_08122_),
    .B1(_08127_),
    .X(_08130_));
 sky130_fd_sc_hd__nand3_1 _18561_ (.A(_08124_),
    .B(_08126_),
    .C(_08127_),
    .Y(_08131_));
 sky130_fd_sc_hd__o21ai_1 _18562_ (.A1(_08123_),
    .A2(_08125_),
    .B1(_08128_),
    .Y(_08132_));
 sky130_fd_sc_hd__o21ai_1 _18563_ (.A1(_08123_),
    .A2(_08125_),
    .B1(_08127_),
    .Y(_08133_));
 sky130_fd_sc_hd__nand3_1 _18564_ (.A(_08124_),
    .B(_08126_),
    .C(_08128_),
    .Y(_08134_));
 sky130_fd_sc_hd__nand3_2 _18565_ (.A(_08133_),
    .B(_08134_),
    .C(net280),
    .Y(_08135_));
 sky130_fd_sc_hd__a311o_2 _18566_ (.A1(_08116_),
    .A2(_08117_),
    .A3(net309),
    .B1(_08119_),
    .C1(net280),
    .X(_08136_));
 sky130_fd_sc_hd__a211o_1 _18567_ (.A1(_08120_),
    .A2(_08121_),
    .B1(net306),
    .C1(net303),
    .X(_08137_));
 sky130_fd_sc_hd__nand3_2 _18568_ (.A(_08132_),
    .B(net280),
    .C(_08131_),
    .Y(_08138_));
 sky130_fd_sc_hd__o221a_2 _18569_ (.A1(_03986_),
    .A2(_03997_),
    .B1(_08122_),
    .B2(net280),
    .C1(_08135_),
    .X(_08139_));
 sky130_fd_sc_hd__a211o_1 _18570_ (.A1(_08137_),
    .A2(_08138_),
    .B1(_04008_),
    .C1(net300),
    .X(_08141_));
 sky130_fd_sc_hd__a21oi_1 _18571_ (.A1(_08135_),
    .A2(_08136_),
    .B1(net319),
    .Y(_08142_));
 sky130_fd_sc_hd__nand3_4 _18572_ (.A(_08138_),
    .B(net320),
    .C(_08137_),
    .Y(_08143_));
 sky130_fd_sc_hd__nand3_4 _18573_ (.A(net319),
    .B(_08135_),
    .C(_08136_),
    .Y(_08144_));
 sky130_fd_sc_hd__a21oi_1 _18574_ (.A1(net325),
    .A2(_07760_),
    .B1(_07763_),
    .Y(_08145_));
 sky130_fd_sc_hd__a22oi_2 _18575_ (.A1(_07422_),
    .A2(_07437_),
    .B1(_07764_),
    .B2(_07747_),
    .Y(_08146_));
 sky130_fd_sc_hd__a21oi_1 _18576_ (.A1(_07763_),
    .A2(_07766_),
    .B1(_07768_),
    .Y(_08147_));
 sky130_fd_sc_hd__o2bb2ai_2 _18577_ (.A1_N(_08143_),
    .A2_N(_08144_),
    .B1(_08145_),
    .B2(_07765_),
    .Y(_08148_));
 sky130_fd_sc_hd__o211ai_4 _18578_ (.A1(_07768_),
    .A2(_08146_),
    .B1(_08144_),
    .C1(_08143_),
    .Y(_08149_));
 sky130_fd_sc_hd__and3_1 _18579_ (.A(_08148_),
    .B(_08149_),
    .C(net275),
    .X(_08150_));
 sky130_fd_sc_hd__nand3_1 _18580_ (.A(_08148_),
    .B(_08149_),
    .C(net275),
    .Y(_08152_));
 sky130_fd_sc_hd__a31o_2 _18581_ (.A1(_08148_),
    .A2(_08149_),
    .A3(net275),
    .B1(_08139_),
    .X(_08153_));
 sky130_fd_sc_hd__and3_1 _18582_ (.A(_05234_),
    .B(_08141_),
    .C(_08152_),
    .X(_08154_));
 sky130_fd_sc_hd__a31oi_4 _18583_ (.A1(net330),
    .A2(_07761_),
    .A3(_07775_),
    .B1(_07784_),
    .Y(_08155_));
 sky130_fd_sc_hd__o21a_1 _18584_ (.A1(_07442_),
    .A2(_07449_),
    .B1(_07780_),
    .X(_08156_));
 sky130_fd_sc_hd__a311oi_4 _18585_ (.A1(_08148_),
    .A2(_08149_),
    .A3(net276),
    .B1(_08139_),
    .C1(net325),
    .Y(_08157_));
 sky130_fd_sc_hd__a311o_2 _18586_ (.A1(_08148_),
    .A2(_08149_),
    .A3(net275),
    .B1(_08139_),
    .C1(net326),
    .X(_08158_));
 sky130_fd_sc_hd__a2bb2oi_2 _18587_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_08141_),
    .B2(_08152_),
    .Y(_08159_));
 sky130_fd_sc_hd__o21ai_4 _18588_ (.A1(_12845_),
    .A2(_12856_),
    .B1(_08153_),
    .Y(_08160_));
 sky130_fd_sc_hd__o211ai_2 _18589_ (.A1(_07779_),
    .A2(_08155_),
    .B1(_08158_),
    .C1(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__o22ai_2 _18590_ (.A1(_07781_),
    .A2(_08156_),
    .B1(_08157_),
    .B2(_08159_),
    .Y(_08163_));
 sky130_fd_sc_hd__nand3_1 _18591_ (.A(_08161_),
    .B(_08163_),
    .C(_05233_),
    .Y(_08164_));
 sky130_fd_sc_hd__o22a_1 _18592_ (.A1(_05228_),
    .A2(_05230_),
    .B1(_08139_),
    .B2(_08150_),
    .X(_08165_));
 sky130_fd_sc_hd__a211o_1 _18593_ (.A1(_08141_),
    .A2(_08152_),
    .B1(net297),
    .C1(_05232_),
    .X(_08166_));
 sky130_fd_sc_hd__o211ai_4 _18594_ (.A1(_07781_),
    .A2(_08156_),
    .B1(_08158_),
    .C1(_08160_),
    .Y(_08167_));
 sky130_fd_sc_hd__o22ai_4 _18595_ (.A1(_07779_),
    .A2(_08155_),
    .B1(_08157_),
    .B2(_08159_),
    .Y(_08168_));
 sky130_fd_sc_hd__nand3_1 _18596_ (.A(_08167_),
    .B(_08168_),
    .C(_05233_),
    .Y(_08169_));
 sky130_fd_sc_hd__a31o_1 _18597_ (.A1(_08167_),
    .A2(_08168_),
    .A3(_05233_),
    .B1(_08165_),
    .X(_08170_));
 sky130_fd_sc_hd__a311oi_2 _18598_ (.A1(_08161_),
    .A2(_08163_),
    .A3(_05233_),
    .B1(_08154_),
    .C1(net331),
    .Y(_08171_));
 sky130_fd_sc_hd__o211ai_4 _18599_ (.A1(_08153_),
    .A2(_05233_),
    .B1(net330),
    .C1(_08164_),
    .Y(_08172_));
 sky130_fd_sc_hd__a311oi_4 _18600_ (.A1(_08167_),
    .A2(_08168_),
    .A3(_05233_),
    .B1(_08165_),
    .C1(net330),
    .Y(_08174_));
 sky130_fd_sc_hd__o211ai_4 _18601_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_08166_),
    .C1(_08169_),
    .Y(_08175_));
 sky130_fd_sc_hd__o21a_1 _18602_ (.A1(_10015_),
    .A2(_07791_),
    .B1(_07798_),
    .X(_08176_));
 sky130_fd_sc_hd__a31o_1 _18603_ (.A1(_09982_),
    .A2(_10004_),
    .A3(_07792_),
    .B1(_07799_),
    .X(_08177_));
 sky130_fd_sc_hd__a21oi_1 _18604_ (.A1(_07797_),
    .A2(_07799_),
    .B1(_07794_),
    .Y(_08178_));
 sky130_fd_sc_hd__o2111ai_4 _18605_ (.A1(_07796_),
    .A2(_07798_),
    .B1(_08172_),
    .C1(_08175_),
    .D1(_07795_),
    .Y(_08179_));
 sky130_fd_sc_hd__o22ai_2 _18606_ (.A1(_07794_),
    .A2(_07806_),
    .B1(_08171_),
    .B2(_08174_),
    .Y(_08180_));
 sky130_fd_sc_hd__o211ai_4 _18607_ (.A1(_05481_),
    .A2(net269),
    .B1(_08179_),
    .C1(_08180_),
    .Y(_08181_));
 sky130_fd_sc_hd__a311o_2 _18608_ (.A1(_08161_),
    .A2(_08163_),
    .A3(_05233_),
    .B1(net246),
    .C1(_08154_),
    .X(_08182_));
 sky130_fd_sc_hd__o2bb2ai_1 _18609_ (.A1_N(_08172_),
    .A2_N(_08175_),
    .B1(_08176_),
    .B2(_07796_),
    .Y(_08183_));
 sky130_fd_sc_hd__o211ai_1 _18610_ (.A1(_07794_),
    .A2(_07806_),
    .B1(_08172_),
    .C1(_08175_),
    .Y(_08185_));
 sky130_fd_sc_hd__nand3_2 _18611_ (.A(_08183_),
    .B(_08185_),
    .C(net246),
    .Y(_08186_));
 sky130_fd_sc_hd__and3_1 _18612_ (.A(_05754_),
    .B(_08182_),
    .C(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__inv_2 _18613_ (.A(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__a2bb2oi_1 _18614_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_08182_),
    .B2(_08186_),
    .Y(_08189_));
 sky130_fd_sc_hd__o211ai_4 _18615_ (.A1(_05485_),
    .A2(_08170_),
    .B1(_08181_),
    .C1(net348),
    .Y(_08190_));
 sky130_fd_sc_hd__o211a_1 _18616_ (.A1(net365),
    .A2(net364),
    .B1(_08182_),
    .C1(_08186_),
    .X(_08191_));
 sky130_fd_sc_hd__o211ai_4 _18617_ (.A1(net365),
    .A2(net364),
    .B1(_08182_),
    .C1(_08186_),
    .Y(_08192_));
 sky130_fd_sc_hd__a22oi_2 _18618_ (.A1(_07478_),
    .A2(_07486_),
    .B1(_07809_),
    .B2(_08907_),
    .Y(_08193_));
 sky130_fd_sc_hd__a21oi_2 _18619_ (.A1(_07813_),
    .A2(_07815_),
    .B1(_07816_),
    .Y(_08194_));
 sky130_fd_sc_hd__o21ai_1 _18620_ (.A1(_08189_),
    .A2(_08191_),
    .B1(_08194_),
    .Y(_08196_));
 sky130_fd_sc_hd__o21ai_1 _18621_ (.A1(_07816_),
    .A2(_08193_),
    .B1(_08192_),
    .Y(_08197_));
 sky130_fd_sc_hd__o211ai_2 _18622_ (.A1(_07816_),
    .A2(_08193_),
    .B1(_08192_),
    .C1(_08190_),
    .Y(_08198_));
 sky130_fd_sc_hd__nand3_2 _18623_ (.A(_08194_),
    .B(_08192_),
    .C(_08190_),
    .Y(_08199_));
 sky130_fd_sc_hd__a21o_1 _18624_ (.A1(_08190_),
    .A2(_08192_),
    .B1(_08194_),
    .X(_08200_));
 sky130_fd_sc_hd__o211ai_2 _18625_ (.A1(net266),
    .A2(_05751_),
    .B1(_08199_),
    .C1(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__o211a_1 _18626_ (.A1(_05485_),
    .A2(_08170_),
    .B1(_08181_),
    .C1(_05754_),
    .X(_08202_));
 sky130_fd_sc_hd__nand3_1 _18627_ (.A(_08196_),
    .B(_08198_),
    .C(net241),
    .Y(_08203_));
 sky130_fd_sc_hd__a31o_2 _18628_ (.A1(_08200_),
    .A2(net241),
    .A3(_08199_),
    .B1(_08187_),
    .X(_08204_));
 sky130_fd_sc_hd__and3_1 _18629_ (.A(_08201_),
    .B(_05995_),
    .C(_08188_),
    .X(_08205_));
 sky130_fd_sc_hd__a311o_1 _18630_ (.A1(_08200_),
    .A2(net241),
    .A3(_08199_),
    .B1(net240),
    .C1(_08187_),
    .X(_08207_));
 sky130_fd_sc_hd__a31oi_4 _18631_ (.A1(_07812_),
    .A2(_07824_),
    .A3(_07888_),
    .B1(_07831_),
    .Y(_08208_));
 sky130_fd_sc_hd__o21a_1 _18632_ (.A1(_07888_),
    .A2(_07825_),
    .B1(_07831_),
    .X(_08209_));
 sky130_fd_sc_hd__a311oi_2 _18633_ (.A1(_08196_),
    .A2(_08198_),
    .A3(net241),
    .B1(_08202_),
    .C1(_08918_),
    .Y(_08210_));
 sky130_fd_sc_hd__nand3b_2 _18634_ (.A_N(_08202_),
    .B(_08203_),
    .C(_08907_),
    .Y(_08211_));
 sky130_fd_sc_hd__a311oi_1 _18635_ (.A1(_08200_),
    .A2(net241),
    .A3(_08199_),
    .B1(_08187_),
    .C1(_08907_),
    .Y(_08212_));
 sky130_fd_sc_hd__o211ai_4 _18636_ (.A1(_08819_),
    .A2(_08841_),
    .B1(_08188_),
    .C1(_08201_),
    .Y(_08213_));
 sky130_fd_sc_hd__o211ai_2 _18637_ (.A1(_07828_),
    .A2(_08208_),
    .B1(_08211_),
    .C1(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__o22ai_2 _18638_ (.A1(_07827_),
    .A2(_08209_),
    .B1(_08210_),
    .B2(_08212_),
    .Y(_08215_));
 sky130_fd_sc_hd__and3_1 _18639_ (.A(net240),
    .B(_08214_),
    .C(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__o211ai_4 _18640_ (.A1(net259),
    .A2(net256),
    .B1(_08214_),
    .C1(_08215_),
    .Y(_08218_));
 sky130_fd_sc_hd__o31a_2 _18641_ (.A1(net259),
    .A2(net256),
    .A3(_08204_),
    .B1(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__or4_1 _18642_ (.A(_06291_),
    .B(_06292_),
    .C(_08205_),
    .D(_08216_),
    .X(_08220_));
 sky130_fd_sc_hd__a21oi_2 _18643_ (.A1(_07842_),
    .A2(_07845_),
    .B1(_07846_),
    .Y(_08221_));
 sky130_fd_sc_hd__o221a_2 _18644_ (.A1(_07844_),
    .A2(_07866_),
    .B1(net240),
    .B2(_08204_),
    .C1(_08218_),
    .X(_08222_));
 sky130_fd_sc_hd__o221ai_4 _18645_ (.A1(_07844_),
    .A2(_07866_),
    .B1(_05996_),
    .B2(_08204_),
    .C1(_08218_),
    .Y(_08223_));
 sky130_fd_sc_hd__a21oi_4 _18646_ (.A1(_08207_),
    .A2(_08218_),
    .B1(_07888_),
    .Y(_08224_));
 sky130_fd_sc_hd__a22o_1 _18647_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_08207_),
    .B2(_08218_),
    .X(_08225_));
 sky130_fd_sc_hd__o2111ai_1 _18648_ (.A1(_07841_),
    .A2(_07843_),
    .B1(_07847_),
    .C1(_08223_),
    .D1(_08225_),
    .Y(_08226_));
 sky130_fd_sc_hd__o21bai_1 _18649_ (.A1(_08222_),
    .A2(_08224_),
    .B1_N(_08221_),
    .Y(_08227_));
 sky130_fd_sc_hd__o211ai_1 _18650_ (.A1(_06291_),
    .A2(_06292_),
    .B1(_08226_),
    .C1(_08227_),
    .Y(_08229_));
 sky130_fd_sc_hd__or3_1 _18651_ (.A(_06291_),
    .B(_06292_),
    .C(_08219_),
    .X(_08230_));
 sky130_fd_sc_hd__o311a_2 _18652_ (.A1(_07503_),
    .A2(_07509_),
    .A3(_07846_),
    .B1(_08223_),
    .C1(_07845_),
    .X(_08231_));
 sky130_fd_sc_hd__nand3b_1 _18653_ (.A_N(_08221_),
    .B(_08223_),
    .C(_08225_),
    .Y(_08232_));
 sky130_fd_sc_hd__o21ai_1 _18654_ (.A1(_08222_),
    .A2(_08224_),
    .B1(_08221_),
    .Y(_08233_));
 sky130_fd_sc_hd__nand3_2 _18655_ (.A(_08233_),
    .B(net212),
    .C(_08232_),
    .Y(_08234_));
 sky130_fd_sc_hd__o31a_2 _18656_ (.A1(_06291_),
    .A2(_06292_),
    .A3(_08219_),
    .B1(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__o221ai_4 _18657_ (.A1(_06989_),
    .A2(net375),
    .B1(net212),
    .B2(_08219_),
    .C1(_08234_),
    .Y(_08236_));
 sky130_fd_sc_hd__o311a_1 _18658_ (.A1(net212),
    .A2(_08205_),
    .A3(_08216_),
    .B1(_08229_),
    .C1(_07044_),
    .X(_08237_));
 sky130_fd_sc_hd__o211ai_1 _18659_ (.A1(_06945_),
    .A2(_06967_),
    .B1(_08220_),
    .C1(_08229_),
    .Y(_08238_));
 sky130_fd_sc_hd__nand3_1 _18660_ (.A(_07925_),
    .B(_08236_),
    .C(_08238_),
    .Y(_08240_));
 sky130_fd_sc_hd__a21o_1 _18661_ (.A1(_08236_),
    .A2(_08238_),
    .B1(_07925_),
    .X(_08241_));
 sky130_fd_sc_hd__o211ai_4 _18662_ (.A1(_06608_),
    .A2(net237),
    .B1(_08240_),
    .C1(_08241_),
    .Y(_08242_));
 sky130_fd_sc_hd__a211o_2 _18663_ (.A1(_08230_),
    .A2(_08234_),
    .B1(_06608_),
    .C1(net237),
    .X(_08243_));
 sky130_fd_sc_hd__o31a_1 _18664_ (.A1(_06608_),
    .A2(net237),
    .A3(_08235_),
    .B1(_08242_),
    .X(_08244_));
 sky130_fd_sc_hd__o311a_1 _18665_ (.A1(_06608_),
    .A2(_08235_),
    .A3(net237),
    .B1(_06904_),
    .C1(_08242_),
    .X(_08245_));
 sky130_fd_sc_hd__o21ai_1 _18666_ (.A1(_06897_),
    .A2(_06898_),
    .B1(_08244_),
    .Y(_08246_));
 sky130_fd_sc_hd__a22oi_4 _18667_ (.A1(_06256_),
    .A2(_06278_),
    .B1(_08242_),
    .B2(_08243_),
    .Y(_08247_));
 sky130_fd_sc_hd__o221a_1 _18668_ (.A1(net381),
    .A2(_06310_),
    .B1(_06612_),
    .B2(_08235_),
    .C1(_08242_),
    .X(_08248_));
 sky130_fd_sc_hd__o221ai_4 _18669_ (.A1(net381),
    .A2(_06310_),
    .B1(_06612_),
    .B2(_08235_),
    .C1(_08242_),
    .Y(_08249_));
 sky130_fd_sc_hd__a21oi_1 _18670_ (.A1(_07873_),
    .A2(_07879_),
    .B1(_07876_),
    .Y(_08251_));
 sky130_fd_sc_hd__a31o_1 _18671_ (.A1(_07870_),
    .A2(_07871_),
    .A3(_07879_),
    .B1(_07876_),
    .X(_08252_));
 sky130_fd_sc_hd__nand3b_1 _18672_ (.A_N(_08247_),
    .B(_08249_),
    .C(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__o21ai_1 _18673_ (.A1(_08247_),
    .A2(_08248_),
    .B1(_08251_),
    .Y(_08254_));
 sky130_fd_sc_hd__o21ai_2 _18674_ (.A1(_08247_),
    .A2(_08248_),
    .B1(_08252_),
    .Y(_08255_));
 sky130_fd_sc_hd__a31oi_4 _18675_ (.A1(_08242_),
    .A2(_08243_),
    .A3(_06332_),
    .B1(_08252_),
    .Y(_08256_));
 sky130_fd_sc_hd__o21ai_2 _18676_ (.A1(_06332_),
    .A2(_08244_),
    .B1(_08256_),
    .Y(_08257_));
 sky130_fd_sc_hd__a22oi_4 _18677_ (.A1(_06900_),
    .A2(_06902_),
    .B1(_08255_),
    .B2(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__o211ai_1 _18678_ (.A1(net230),
    .A2(_06901_),
    .B1(_08253_),
    .C1(_08254_),
    .Y(_08259_));
 sky130_fd_sc_hd__nand3_1 _18679_ (.A(_08255_),
    .B(_08257_),
    .C(net208),
    .Y(_08260_));
 sky130_fd_sc_hd__o211ai_2 _18680_ (.A1(_05556_),
    .A2(_07887_),
    .B1(_07885_),
    .C1(_07883_),
    .Y(_08262_));
 sky130_fd_sc_hd__o31a_1 _18681_ (.A1(_05501_),
    .A2(_05523_),
    .A3(_07886_),
    .B1(_08262_),
    .X(_08263_));
 sky130_fd_sc_hd__a21oi_1 _18682_ (.A1(_07890_),
    .A2(_08262_),
    .B1(_05851_),
    .Y(_08264_));
 sky130_fd_sc_hd__o21ai_1 _18683_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_08263_),
    .Y(_08265_));
 sky130_fd_sc_hd__a31oi_1 _18684_ (.A1(_08262_),
    .A2(_05851_),
    .A3(_07890_),
    .B1(_07232_),
    .Y(_08266_));
 sky130_fd_sc_hd__o21ai_2 _18685_ (.A1(_05851_),
    .A2(_08263_),
    .B1(_08266_),
    .Y(_08267_));
 sky130_fd_sc_hd__o211ai_2 _18686_ (.A1(net208),
    .A2(_08244_),
    .B1(_08260_),
    .C1(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__o31a_1 _18687_ (.A1(_08245_),
    .A2(_08267_),
    .A3(_08258_),
    .B1(_08268_),
    .X(_08269_));
 sky130_fd_sc_hd__o31ai_4 _18688_ (.A1(_08245_),
    .A2(_08267_),
    .A3(_08258_),
    .B1(_08268_),
    .Y(_08270_));
 sky130_fd_sc_hd__a2bb2oi_1 _18689_ (.A1_N(_05447_),
    .A2_N(_05469_),
    .B1(_07897_),
    .B2(_07904_),
    .Y(_08271_));
 sky130_fd_sc_hd__o21ai_4 _18690_ (.A1(_07898_),
    .A2(_07903_),
    .B1(_05556_),
    .Y(_08273_));
 sky130_fd_sc_hd__o221a_1 _18691_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_07541_),
    .B2(_07900_),
    .C1(_07897_),
    .X(_08274_));
 sky130_fd_sc_hd__o221ai_4 _18692_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_07541_),
    .B2(_07900_),
    .C1(_07897_),
    .Y(_08275_));
 sky130_fd_sc_hd__a31oi_1 _18693_ (.A1(_07904_),
    .A2(_05545_),
    .A3(_07897_),
    .B1(_07550_),
    .Y(_08276_));
 sky130_fd_sc_hd__o21ai_1 _18694_ (.A1(_07544_),
    .A2(net184),
    .B1(_08275_),
    .Y(_08277_));
 sky130_fd_sc_hd__a31o_2 _18695_ (.A1(_08273_),
    .A2(_08275_),
    .A3(net163),
    .B1(_08270_),
    .X(_08278_));
 sky130_fd_sc_hd__nand4_4 _18696_ (.A(_08270_),
    .B(_08273_),
    .C(_08275_),
    .D(net163),
    .Y(_08279_));
 sky130_fd_sc_hd__nand3_1 _18697_ (.A(_08269_),
    .B(_08273_),
    .C(_08276_),
    .Y(_08280_));
 sky130_fd_sc_hd__o21ai_1 _18698_ (.A1(_08271_),
    .A2(_08277_),
    .B1(_08270_),
    .Y(_08281_));
 sky130_fd_sc_hd__nand3_4 _18699_ (.A(_08281_),
    .B(_05239_),
    .C(_08280_),
    .Y(_08282_));
 sky130_fd_sc_hd__nand3_2 _18700_ (.A(_05250_),
    .B(_08278_),
    .C(_08279_),
    .Y(_08284_));
 sky130_fd_sc_hd__o21ai_2 _18701_ (.A1(_03289_),
    .A2(_07907_),
    .B1(_08282_),
    .Y(_08285_));
 sky130_fd_sc_hd__o2bb2ai_1 _18702_ (.A1_N(_08282_),
    .A2_N(_08284_),
    .B1(_03289_),
    .B2(_07907_),
    .Y(_08286_));
 sky130_fd_sc_hd__nand4_1 _18703_ (.A(_08284_),
    .B(_07906_),
    .C(net1),
    .D(_08282_),
    .Y(_08287_));
 sky130_fd_sc_hd__o211ai_2 _18704_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_08286_),
    .C1(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__a211o_1 _18705_ (.A1(_08278_),
    .A2(_08279_),
    .B1(_07912_),
    .C1(_07914_),
    .X(_08289_));
 sky130_fd_sc_hd__a21o_2 _18706_ (.A1(_08288_),
    .A2(_08289_),
    .B1(_03289_),
    .X(_08290_));
 sky130_fd_sc_hd__nand3_1 _18707_ (.A(_03289_),
    .B(_08288_),
    .C(_08289_),
    .Y(_08291_));
 sky130_fd_sc_hd__or4_4 _18708_ (.A(net45),
    .B(net46),
    .C(net47),
    .D(_07226_),
    .X(_08292_));
 sky130_fd_sc_hd__and3_2 _18709_ (.A(_08292_),
    .B(net48),
    .C(net409),
    .X(_08293_));
 sky130_fd_sc_hd__a21oi_4 _18710_ (.A1(_08292_),
    .A2(net409),
    .B1(net48),
    .Y(_08295_));
 sky130_fd_sc_hd__a21boi_4 _18711_ (.A1(_08292_),
    .A2(net409),
    .B1_N(net48),
    .Y(_08296_));
 sky130_fd_sc_hd__a21bo_4 _18712_ (.A1(_08292_),
    .A2(net409),
    .B1_N(net48),
    .X(_08297_));
 sky130_fd_sc_hd__and3b_4 _18713_ (.A_N(net48),
    .B(_08292_),
    .C(net409),
    .X(_08298_));
 sky130_fd_sc_hd__nand3b_4 _18714_ (.A_N(net48),
    .B(_08292_),
    .C(net409),
    .Y(_08299_));
 sky130_fd_sc_hd__nand2_8 _18715_ (.A(_08297_),
    .B(_08299_),
    .Y(_08300_));
 sky130_fd_sc_hd__nor2_8 _18716_ (.A(net180),
    .B(_08298_),
    .Y(_08301_));
 sky130_fd_sc_hd__o2bb2a_1 _18717_ (.A1_N(_08290_),
    .A2_N(_08291_),
    .B1(net180),
    .B2(_08298_),
    .X(_08302_));
 sky130_fd_sc_hd__a31o_1 _18718_ (.A1(_08288_),
    .A2(_08289_),
    .A3(_08301_),
    .B1(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__xnor2_1 _18719_ (.A(_07924_),
    .B(_08303_),
    .Y(net80));
 sky130_fd_sc_hd__nor3b_1 _18720_ (.A(_07553_),
    .B(_07920_),
    .C_N(_08303_),
    .Y(_08305_));
 sky130_fd_sc_hd__or4_4 _18721_ (.A(net14),
    .B(net15),
    .C(net16),
    .D(_07240_),
    .X(_08306_));
 sky130_fd_sc_hd__and3b_4 _18722_ (.A_N(net17),
    .B(_08306_),
    .C(net410),
    .X(_08307_));
 sky130_fd_sc_hd__nand3b_4 _18723_ (.A_N(net17),
    .B(_08306_),
    .C(net410),
    .Y(_08308_));
 sky130_fd_sc_hd__a21boi_4 _18724_ (.A1(_08306_),
    .A2(net410),
    .B1_N(net17),
    .Y(_08309_));
 sky130_fd_sc_hd__a21bo_4 _18725_ (.A1(_08306_),
    .A2(net410),
    .B1_N(net17),
    .X(_08310_));
 sky130_fd_sc_hd__o311a_4 _18726_ (.A1(net15),
    .A2(net16),
    .A3(_07554_),
    .B1(net17),
    .C1(net410),
    .X(_08311_));
 sky130_fd_sc_hd__a21oi_4 _18727_ (.A1(_08306_),
    .A2(net410),
    .B1(net17),
    .Y(_08312_));
 sky130_fd_sc_hd__nor2_8 _18728_ (.A(_08307_),
    .B(net216),
    .Y(_08313_));
 sky130_fd_sc_hd__nor2_8 _18729_ (.A(_08311_),
    .B(net215),
    .Y(_08314_));
 sky130_fd_sc_hd__a21oi_2 _18730_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_03178_),
    .Y(_08316_));
 sky130_fd_sc_hd__or3_4 _18731_ (.A(_03178_),
    .B(_08311_),
    .C(_08312_),
    .X(_08317_));
 sky130_fd_sc_hd__or3_1 _18732_ (.A(_07928_),
    .B(_07930_),
    .C(_08316_),
    .X(_08318_));
 sky130_fd_sc_hd__o31a_1 _18733_ (.A1(_07938_),
    .A2(_08311_),
    .A3(_08312_),
    .B1(_08318_),
    .X(_08319_));
 sky130_fd_sc_hd__o21ai_1 _18734_ (.A1(_07938_),
    .A2(net199),
    .B1(_08318_),
    .Y(_08320_));
 sky130_fd_sc_hd__o211ai_2 _18735_ (.A1(_07935_),
    .A2(_07566_),
    .B1(_07569_),
    .C1(_07573_),
    .Y(_08321_));
 sky130_fd_sc_hd__o2bb2ai_1 _18736_ (.A1_N(_07569_),
    .A2_N(_07573_),
    .B1(_07937_),
    .B2(net202),
    .Y(_08322_));
 sky130_fd_sc_hd__o211ai_2 _18737_ (.A1(_07566_),
    .A2(_07935_),
    .B1(_08320_),
    .C1(_08322_),
    .Y(_08323_));
 sky130_fd_sc_hd__o211ai_4 _18738_ (.A1(net202),
    .A2(_07937_),
    .B1(_08319_),
    .C1(_08321_),
    .Y(_08324_));
 sky130_fd_sc_hd__o32a_2 _18739_ (.A1(_03178_),
    .A2(_08311_),
    .A3(_08312_),
    .B1(_05130_),
    .B2(_05152_),
    .X(_08325_));
 sky130_fd_sc_hd__a22o_1 _18740_ (.A1(_05141_),
    .A2(_05163_),
    .B1(net198),
    .B2(net33),
    .X(_08327_));
 sky130_fd_sc_hd__a21oi_4 _18741_ (.A1(_08323_),
    .A2(_08324_),
    .B1(_05185_),
    .Y(_08328_));
 sky130_fd_sc_hd__a2111oi_4 _18742_ (.A1(_05185_),
    .A2(_08317_),
    .B1(_08328_),
    .C1(_05348_),
    .D1(net401),
    .Y(_08329_));
 sky130_fd_sc_hd__o21ai_2 _18743_ (.A1(_08325_),
    .A2(_08328_),
    .B1(_07564_),
    .Y(_08330_));
 sky130_fd_sc_hd__a21oi_1 _18744_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_08328_),
    .Y(_08331_));
 sky130_fd_sc_hd__or3_1 _18745_ (.A(_07560_),
    .B(_07562_),
    .C(_08328_),
    .X(_08332_));
 sky130_fd_sc_hd__a221o_2 _18746_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_08317_),
    .B2(_05185_),
    .C1(_08328_),
    .X(_08333_));
 sky130_fd_sc_hd__nand2_4 _18747_ (.A(_08330_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__a22oi_4 _18748_ (.A1(_07950_),
    .A2(_07940_),
    .B1(_07957_),
    .B2(_07954_),
    .Y(_08335_));
 sky130_fd_sc_hd__o2bb2ai_1 _18749_ (.A1_N(_07954_),
    .A2_N(_07957_),
    .B1(_07939_),
    .B2(_07951_),
    .Y(_08336_));
 sky130_fd_sc_hd__o311a_1 _18750_ (.A1(net224),
    .A2(_07939_),
    .A3(_07946_),
    .B1(_07958_),
    .C1(_08334_),
    .X(_08338_));
 sky130_fd_sc_hd__o211ai_2 _18751_ (.A1(_07951_),
    .A2(_07939_),
    .B1(_08334_),
    .C1(_07958_),
    .Y(_08339_));
 sky130_fd_sc_hd__and3_1 _18752_ (.A(_08330_),
    .B(_08333_),
    .C(_08336_),
    .X(_08340_));
 sky130_fd_sc_hd__o211a_1 _18753_ (.A1(_08334_),
    .A2(_08335_),
    .B1(_08339_),
    .C1(_05403_),
    .X(_08341_));
 sky130_fd_sc_hd__o211ai_2 _18754_ (.A1(_08334_),
    .A2(_08335_),
    .B1(_08339_),
    .C1(_05403_),
    .Y(_08342_));
 sky130_fd_sc_hd__o211a_1 _18755_ (.A1(_08325_),
    .A2(_08328_),
    .B1(_05359_),
    .C1(_05381_),
    .X(_08343_));
 sky130_fd_sc_hd__o22a_1 _18756_ (.A1(_05348_),
    .A2(net401),
    .B1(_08338_),
    .B2(_08340_),
    .X(_08344_));
 sky130_fd_sc_hd__o31a_1 _18757_ (.A1(_05403_),
    .A2(_08325_),
    .A3(_08328_),
    .B1(_08342_),
    .X(_08345_));
 sky130_fd_sc_hd__o22a_1 _18758_ (.A1(_05654_),
    .A2(_05665_),
    .B1(_08329_),
    .B2(_08341_),
    .X(_08346_));
 sky130_fd_sc_hd__or4_4 _18759_ (.A(_05676_),
    .B(_05698_),
    .C(_08343_),
    .D(_08344_),
    .X(_08347_));
 sky130_fd_sc_hd__o22a_1 _18760_ (.A1(_07242_),
    .A2(_07243_),
    .B1(_08329_),
    .B2(_08341_),
    .X(_08349_));
 sky130_fd_sc_hd__o22ai_2 _18761_ (.A1(_07242_),
    .A2(_07243_),
    .B1(_08329_),
    .B2(_08341_),
    .Y(_08350_));
 sky130_fd_sc_hd__o21ai_2 _18762_ (.A1(_07244_),
    .A2(_07245_),
    .B1(_08342_),
    .Y(_08351_));
 sky130_fd_sc_hd__o21a_2 _18763_ (.A1(_08329_),
    .A2(_08351_),
    .B1(_08350_),
    .X(_08352_));
 sky130_fd_sc_hd__o21ai_2 _18764_ (.A1(_08329_),
    .A2(_08351_),
    .B1(_08350_),
    .Y(_08353_));
 sky130_fd_sc_hd__a31oi_1 _18765_ (.A1(_07971_),
    .A2(_07978_),
    .A3(_07980_),
    .B1(_07967_),
    .Y(_08354_));
 sky130_fd_sc_hd__o22ai_4 _18766_ (.A1(net227),
    .A2(_07963_),
    .B1(_07983_),
    .B2(_07977_),
    .Y(_08355_));
 sky130_fd_sc_hd__a21oi_1 _18767_ (.A1(_07968_),
    .A2(_07985_),
    .B1(_08353_),
    .Y(_08356_));
 sky130_fd_sc_hd__nand2_2 _18768_ (.A(_08355_),
    .B(_08352_),
    .Y(_08357_));
 sky130_fd_sc_hd__o221ai_4 _18769_ (.A1(net227),
    .A2(_07963_),
    .B1(_07983_),
    .B2(_07977_),
    .C1(_08353_),
    .Y(_08358_));
 sky130_fd_sc_hd__o221a_1 _18770_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_08352_),
    .B2(_08355_),
    .C1(_08357_),
    .X(_08360_));
 sky130_fd_sc_hd__nand3_1 _18771_ (.A(_08357_),
    .B(_08358_),
    .C(net358),
    .Y(_08361_));
 sky130_fd_sc_hd__a31oi_4 _18772_ (.A1(_08357_),
    .A2(_08358_),
    .A3(net358),
    .B1(_08346_),
    .Y(_08362_));
 sky130_fd_sc_hd__or3_2 _18773_ (.A(_06793_),
    .B(_06815_),
    .C(_08362_),
    .X(_08363_));
 sky130_fd_sc_hd__inv_2 _18774_ (.A(_08363_),
    .Y(_08364_));
 sky130_fd_sc_hd__a2bb2oi_4 _18775_ (.A1_N(_06914_),
    .A2_N(_06916_),
    .B1(_08347_),
    .B2(_08361_),
    .Y(_08365_));
 sky130_fd_sc_hd__o22ai_1 _18776_ (.A1(_06914_),
    .A2(_06916_),
    .B1(_08346_),
    .B2(_08360_),
    .Y(_08366_));
 sky130_fd_sc_hd__a31oi_2 _18777_ (.A1(_08357_),
    .A2(_08358_),
    .A3(net358),
    .B1(net225),
    .Y(_08367_));
 sky130_fd_sc_hd__o221a_1 _18778_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_08345_),
    .B2(net358),
    .C1(_08361_),
    .X(_08368_));
 sky130_fd_sc_hd__a311o_1 _18779_ (.A1(_08357_),
    .A2(_08358_),
    .A3(net358),
    .B1(net225),
    .C1(_08346_),
    .X(_08369_));
 sky130_fd_sc_hd__a21oi_4 _18780_ (.A1(_08347_),
    .A2(_08367_),
    .B1(_08365_),
    .Y(_08371_));
 sky130_fd_sc_hd__o2111ai_2 _18781_ (.A1(_07295_),
    .A2(_07286_),
    .B1(_06971_),
    .C1(_06968_),
    .D1(_07293_),
    .Y(_08372_));
 sky130_fd_sc_hd__nor3_2 _18782_ (.A(_07617_),
    .B(_07621_),
    .C(_08372_),
    .Y(_08373_));
 sky130_fd_sc_hd__nand2_1 _18783_ (.A(_08373_),
    .B(_07998_),
    .Y(_08374_));
 sky130_fd_sc_hd__a41oi_4 _18784_ (.A1(_07998_),
    .A2(_07623_),
    .A3(_07298_),
    .A4(_06972_),
    .B1(_07999_),
    .Y(_08375_));
 sky130_fd_sc_hd__o211a_1 _18785_ (.A1(_07996_),
    .A2(_07994_),
    .B1(_08374_),
    .C1(_08000_),
    .X(_08376_));
 sky130_fd_sc_hd__o211ai_4 _18786_ (.A1(_07996_),
    .A2(_07994_),
    .B1(_08374_),
    .C1(_08000_),
    .Y(_08377_));
 sky130_fd_sc_hd__and4b_1 _18787_ (.A_N(_08372_),
    .B(_07622_),
    .C(_07618_),
    .D(_06987_),
    .X(_08378_));
 sky130_fd_sc_hd__o211ai_2 _18788_ (.A1(_06981_),
    .A2(_06984_),
    .B1(_08373_),
    .C1(_08000_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand4_4 _18789_ (.A(_08373_),
    .B(_08000_),
    .C(_07998_),
    .D(_06987_),
    .Y(_08380_));
 sky130_fd_sc_hd__a22oi_2 _18790_ (.A1(_08001_),
    .A2(_08378_),
    .B1(_08002_),
    .B2(_08375_),
    .Y(_08382_));
 sky130_fd_sc_hd__o2bb2ai_4 _18791_ (.A1_N(_08375_),
    .A2_N(_08002_),
    .B1(_07996_),
    .B2(_08379_),
    .Y(_08383_));
 sky130_fd_sc_hd__nand3_1 _18792_ (.A(_08366_),
    .B(_08369_),
    .C(_08380_),
    .Y(_08384_));
 sky130_fd_sc_hd__nand3_4 _18793_ (.A(_08371_),
    .B(_08377_),
    .C(_08380_),
    .Y(_08385_));
 sky130_fd_sc_hd__o21ai_1 _18794_ (.A1(_08365_),
    .A2(_08368_),
    .B1(_08383_),
    .Y(_08386_));
 sky130_fd_sc_hd__o221a_1 _18795_ (.A1(net379),
    .A2(net378),
    .B1(_08371_),
    .B2(_08382_),
    .C1(_08385_),
    .X(_08387_));
 sky130_fd_sc_hd__o221ai_4 _18796_ (.A1(net379),
    .A2(net378),
    .B1(_08371_),
    .B2(_08382_),
    .C1(_08385_),
    .Y(_08388_));
 sky130_fd_sc_hd__o31a_1 _18797_ (.A1(_06793_),
    .A2(_06815_),
    .A3(_08362_),
    .B1(_08388_),
    .X(_08389_));
 sky130_fd_sc_hd__inv_2 _18798_ (.A(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__a211o_2 _18799_ (.A1(_08363_),
    .A2(_08388_),
    .B1(_07691_),
    .C1(net371),
    .X(_08391_));
 sky130_fd_sc_hd__inv_2 _18800_ (.A(_08391_),
    .Y(_08393_));
 sky130_fd_sc_hd__o211a_1 _18801_ (.A1(_07641_),
    .A2(_07638_),
    .B1(_07637_),
    .C1(_08009_),
    .X(_08394_));
 sky130_fd_sc_hd__nand2_1 _18802_ (.A(_08014_),
    .B(_08009_),
    .Y(_08395_));
 sky130_fd_sc_hd__o32ai_4 _18803_ (.A1(net251),
    .A2(_07991_),
    .A3(_08004_),
    .B1(_08007_),
    .B2(_08015_),
    .Y(_08396_));
 sky130_fd_sc_hd__a31oi_1 _18804_ (.A1(_08386_),
    .A2(net357),
    .A3(_08385_),
    .B1(net232),
    .Y(_08397_));
 sky130_fd_sc_hd__o211a_2 _18805_ (.A1(net357),
    .A2(_08362_),
    .B1(net234),
    .C1(_08388_),
    .X(_08398_));
 sky130_fd_sc_hd__o211ai_4 _18806_ (.A1(net357),
    .A2(_08362_),
    .B1(net234),
    .C1(_08388_),
    .Y(_08399_));
 sky130_fd_sc_hd__a2bb2oi_2 _18807_ (.A1_N(_06622_),
    .A2_N(_06624_),
    .B1(_08363_),
    .B2(_08388_),
    .Y(_08400_));
 sky130_fd_sc_hd__o22ai_4 _18808_ (.A1(_06622_),
    .A2(_06624_),
    .B1(_08364_),
    .B2(_08387_),
    .Y(_08401_));
 sky130_fd_sc_hd__a211oi_1 _18809_ (.A1(_08397_),
    .A2(_08363_),
    .B1(_08396_),
    .C1(_08400_),
    .Y(_08402_));
 sky130_fd_sc_hd__o2111ai_4 _18810_ (.A1(net251),
    .A2(_08006_),
    .B1(_08395_),
    .C1(_08399_),
    .D1(_08401_),
    .Y(_08404_));
 sky130_fd_sc_hd__a22oi_1 _18811_ (.A1(_08012_),
    .A2(_08395_),
    .B1(_08399_),
    .B2(_08401_),
    .Y(_08405_));
 sky130_fd_sc_hd__o22ai_2 _18812_ (.A1(_08011_),
    .A2(_08394_),
    .B1(_08398_),
    .B2(_08400_),
    .Y(_08406_));
 sky130_fd_sc_hd__nand3_2 _18813_ (.A(_08406_),
    .B(net355),
    .C(_08404_),
    .Y(_08407_));
 sky130_fd_sc_hd__o22ai_1 _18814_ (.A1(_07691_),
    .A2(net371),
    .B1(_08402_),
    .B2(_08405_),
    .Y(_08408_));
 sky130_fd_sc_hd__o31a_1 _18815_ (.A1(_07691_),
    .A2(net371),
    .A3(_08389_),
    .B1(_08407_),
    .X(_08409_));
 sky130_fd_sc_hd__inv_2 _18816_ (.A(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__a2bb2oi_4 _18817_ (.A1_N(_06305_),
    .A2_N(net283),
    .B1(_08391_),
    .B2(_08407_),
    .Y(_08411_));
 sky130_fd_sc_hd__o211ai_2 _18818_ (.A1(_08390_),
    .A2(net355),
    .B1(net251),
    .C1(_08408_),
    .Y(_08412_));
 sky130_fd_sc_hd__a31oi_1 _18819_ (.A1(_08404_),
    .A2(_08406_),
    .A3(net355),
    .B1(net251),
    .Y(_08413_));
 sky130_fd_sc_hd__a31o_1 _18820_ (.A1(_08406_),
    .A2(net355),
    .A3(_08404_),
    .B1(net251),
    .X(_08415_));
 sky130_fd_sc_hd__o211a_1 _18821_ (.A1(net355),
    .A2(_08389_),
    .B1(_06314_),
    .C1(_08407_),
    .X(_08416_));
 sky130_fd_sc_hd__nand3_2 _18822_ (.A(_08407_),
    .B(_06314_),
    .C(_08391_),
    .Y(_08417_));
 sky130_fd_sc_hd__a21oi_1 _18823_ (.A1(_08391_),
    .A2(_08413_),
    .B1(_08411_),
    .Y(_08418_));
 sky130_fd_sc_hd__o211ai_4 _18824_ (.A1(_08032_),
    .A2(_07662_),
    .B1(_07654_),
    .C1(_08027_),
    .Y(_08419_));
 sky130_fd_sc_hd__o22a_1 _18825_ (.A1(_08028_),
    .A2(_08022_),
    .B1(_08026_),
    .B2(_08033_),
    .X(_08420_));
 sky130_fd_sc_hd__o21ai_1 _18826_ (.A1(net253),
    .A2(_08025_),
    .B1(_08419_),
    .Y(_08421_));
 sky130_fd_sc_hd__o211ai_1 _18827_ (.A1(_08415_),
    .A2(_08393_),
    .B1(_08412_),
    .C1(_08421_),
    .Y(_08422_));
 sky130_fd_sc_hd__o21ai_1 _18828_ (.A1(_08411_),
    .A2(_08416_),
    .B1(_08420_),
    .Y(_08423_));
 sky130_fd_sc_hd__nand3_1 _18829_ (.A(_08423_),
    .B(net338),
    .C(_08422_),
    .Y(_08424_));
 sky130_fd_sc_hd__a211o_1 _18830_ (.A1(_08391_),
    .A2(_08407_),
    .B1(net353),
    .C1(net352),
    .X(_08426_));
 sky130_fd_sc_hd__o21ai_1 _18831_ (.A1(_08411_),
    .A2(_08416_),
    .B1(_08421_),
    .Y(_08427_));
 sky130_fd_sc_hd__nand4_1 _18832_ (.A(_08031_),
    .B(_08412_),
    .C(_08417_),
    .D(_08419_),
    .Y(_08428_));
 sky130_fd_sc_hd__nand3_2 _18833_ (.A(_08427_),
    .B(_08428_),
    .C(net338),
    .Y(_08429_));
 sky130_fd_sc_hd__o21ai_1 _18834_ (.A1(net338),
    .A2(_08409_),
    .B1(_08429_),
    .Y(_08430_));
 sky130_fd_sc_hd__o31a_4 _18835_ (.A1(net353),
    .A2(net352),
    .A3(_08409_),
    .B1(_08429_),
    .X(_08431_));
 sky130_fd_sc_hd__o211ai_4 _18836_ (.A1(_08410_),
    .A2(net338),
    .B1(net253),
    .C1(_08424_),
    .Y(_08432_));
 sky130_fd_sc_hd__nand3_4 _18837_ (.A(_08429_),
    .B(net254),
    .C(_08426_),
    .Y(_08433_));
 sky130_fd_sc_hd__nand2_2 _18838_ (.A(_08432_),
    .B(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__o2bb2ai_2 _18839_ (.A1_N(_08054_),
    .A2_N(_08056_),
    .B1(net262),
    .B2(_08042_),
    .Y(_08435_));
 sky130_fd_sc_hd__a31oi_2 _18840_ (.A1(_08047_),
    .A2(_08054_),
    .A3(_08056_),
    .B1(_08044_),
    .Y(_08437_));
 sky130_fd_sc_hd__o311a_2 _18841_ (.A1(_05765_),
    .A2(net289),
    .A3(_08042_),
    .B1(_08060_),
    .C1(_08434_),
    .X(_08438_));
 sky130_fd_sc_hd__o211ai_2 _18842_ (.A1(net262),
    .A2(_08042_),
    .B1(_08060_),
    .C1(_08434_),
    .Y(_08439_));
 sky130_fd_sc_hd__o2111ai_2 _18843_ (.A1(net261),
    .A2(_08043_),
    .B1(_08432_),
    .C1(_08433_),
    .D1(_08435_),
    .Y(_08440_));
 sky130_fd_sc_hd__o21ai_4 _18844_ (.A1(_08434_),
    .A2(_08437_),
    .B1(net336),
    .Y(_08441_));
 sky130_fd_sc_hd__nand3_2 _18845_ (.A(_08440_),
    .B(net336),
    .C(_08439_),
    .Y(_08442_));
 sky130_fd_sc_hd__or3_2 _18846_ (.A(_09785_),
    .B(net349),
    .C(_08431_),
    .X(_08443_));
 sky130_fd_sc_hd__o22ai_4 _18847_ (.A1(net336),
    .A2(_08431_),
    .B1(_08438_),
    .B2(_08441_),
    .Y(_08444_));
 sky130_fd_sc_hd__inv_2 _18848_ (.A(_08444_),
    .Y(_08445_));
 sky130_fd_sc_hd__o2111ai_2 _18849_ (.A1(_07060_),
    .A2(_07050_),
    .B1(_07059_),
    .C1(_07359_),
    .D1(_07363_),
    .Y(_08446_));
 sky130_fd_sc_hd__a211oi_1 _18850_ (.A1(_07675_),
    .A2(_07694_),
    .B1(_08446_),
    .C1(_07697_),
    .Y(_08448_));
 sky130_fd_sc_hd__nand2_1 _18851_ (.A(_08073_),
    .B(_08448_),
    .Y(_08449_));
 sky130_fd_sc_hd__o211ai_4 _18852_ (.A1(_08078_),
    .A2(_08072_),
    .B1(_08076_),
    .C1(_08449_),
    .Y(_08450_));
 sky130_fd_sc_hd__and4b_1 _18853_ (.A_N(_08446_),
    .B(_07698_),
    .C(_07696_),
    .D(_07072_),
    .X(_08451_));
 sky130_fd_sc_hd__o211ai_2 _18854_ (.A1(net267),
    .A2(_08067_),
    .B1(_08448_),
    .C1(_07072_),
    .Y(_08452_));
 sky130_fd_sc_hd__nand3_4 _18855_ (.A(_08451_),
    .B(_08076_),
    .C(_08073_),
    .Y(_08453_));
 sky130_fd_sc_hd__o21ai_4 _18856_ (.A1(_08072_),
    .A2(_08452_),
    .B1(_08450_),
    .Y(_08454_));
 sky130_fd_sc_hd__inv_2 _18857_ (.A(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__a22oi_4 _18858_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_08442_),
    .B2(_08443_),
    .Y(_08456_));
 sky130_fd_sc_hd__o21ai_2 _18859_ (.A1(_05760_),
    .A2(net290),
    .B1(_08444_),
    .Y(_08457_));
 sky130_fd_sc_hd__a31oi_1 _18860_ (.A1(_08439_),
    .A2(_08440_),
    .A3(net336),
    .B1(net261),
    .Y(_08459_));
 sky130_fd_sc_hd__o221a_1 _18861_ (.A1(net336),
    .A2(_08431_),
    .B1(_08438_),
    .B2(_08441_),
    .C1(net262),
    .X(_08460_));
 sky130_fd_sc_hd__o221ai_4 _18862_ (.A1(net336),
    .A2(_08431_),
    .B1(_08438_),
    .B2(_08441_),
    .C1(net262),
    .Y(_08461_));
 sky130_fd_sc_hd__a21oi_2 _18863_ (.A1(_08443_),
    .A2(_08459_),
    .B1(_08456_),
    .Y(_08462_));
 sky130_fd_sc_hd__nand2_1 _18864_ (.A(_08457_),
    .B(_08461_),
    .Y(_08463_));
 sky130_fd_sc_hd__a21oi_2 _18865_ (.A1(_08450_),
    .A2(_08453_),
    .B1(_08463_),
    .Y(_08464_));
 sky130_fd_sc_hd__o22ai_4 _18866_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_08462_),
    .B2(_08454_),
    .Y(_08465_));
 sky130_fd_sc_hd__o2bb2ai_2 _18867_ (.A1_N(_08450_),
    .A2_N(_08453_),
    .B1(_08456_),
    .B2(_08460_),
    .Y(_08466_));
 sky130_fd_sc_hd__nand4_4 _18868_ (.A(_08450_),
    .B(_08453_),
    .C(_08457_),
    .D(_08461_),
    .Y(_08467_));
 sky130_fd_sc_hd__nand3_1 _18869_ (.A(_08466_),
    .B(_08467_),
    .C(net333),
    .Y(_08468_));
 sky130_fd_sc_hd__a21oi_1 _18870_ (.A1(_08442_),
    .A2(_08443_),
    .B1(net333),
    .Y(_08470_));
 sky130_fd_sc_hd__a211o_1 _18871_ (.A1(_08442_),
    .A2(_08443_),
    .B1(_11046_),
    .C1(_11057_),
    .X(_08471_));
 sky130_fd_sc_hd__o221a_4 _18872_ (.A1(net333),
    .A2(_08444_),
    .B1(_08464_),
    .B2(_08465_),
    .C1(_12703_),
    .X(_08472_));
 sky130_fd_sc_hd__a211o_2 _18873_ (.A1(_08468_),
    .A2(_08471_),
    .B1(_12670_),
    .C1(_12681_),
    .X(_08473_));
 sky130_fd_sc_hd__a311oi_4 _18874_ (.A1(_08466_),
    .A2(_08467_),
    .A3(net333),
    .B1(_08470_),
    .C1(net291),
    .Y(_08474_));
 sky130_fd_sc_hd__nand3_4 _18875_ (.A(_08468_),
    .B(_08471_),
    .C(net267),
    .Y(_08475_));
 sky130_fd_sc_hd__o221a_1 _18876_ (.A1(net333),
    .A2(_08444_),
    .B1(_08464_),
    .B2(_08465_),
    .C1(net291),
    .X(_08476_));
 sky130_fd_sc_hd__o221ai_4 _18877_ (.A1(net333),
    .A2(_08444_),
    .B1(_08464_),
    .B2(_08465_),
    .C1(net291),
    .Y(_08477_));
 sky130_fd_sc_hd__o22a_1 _18878_ (.A1(net295),
    .A2(_08086_),
    .B1(_08088_),
    .B2(_07708_),
    .X(_08478_));
 sky130_fd_sc_hd__o32a_1 _18879_ (.A1(_05242_),
    .A2(net314),
    .A3(_08087_),
    .B1(_08090_),
    .B2(_08094_),
    .X(_08479_));
 sky130_fd_sc_hd__a21oi_2 _18880_ (.A1(_08090_),
    .A2(_08093_),
    .B1(_08094_),
    .Y(_08481_));
 sky130_fd_sc_hd__o2bb2ai_4 _18881_ (.A1_N(_08475_),
    .A2_N(_08477_),
    .B1(_08478_),
    .B2(_08092_),
    .Y(_08482_));
 sky130_fd_sc_hd__nand3_4 _18882_ (.A(_08479_),
    .B(_08477_),
    .C(_08475_),
    .Y(_08483_));
 sky130_fd_sc_hd__o311a_1 _18883_ (.A1(_08474_),
    .A2(_08481_),
    .A3(_08476_),
    .B1(net312),
    .C1(_08482_),
    .X(_08484_));
 sky130_fd_sc_hd__nand3_1 _18884_ (.A(_08482_),
    .B(_08483_),
    .C(net312),
    .Y(_08485_));
 sky130_fd_sc_hd__a31oi_4 _18885_ (.A1(_08482_),
    .A2(_08483_),
    .A3(net312),
    .B1(_08472_),
    .Y(_08486_));
 sky130_fd_sc_hd__a31o_1 _18886_ (.A1(_08482_),
    .A2(_08483_),
    .A3(net312),
    .B1(_08472_),
    .X(_08487_));
 sky130_fd_sc_hd__o221a_1 _18887_ (.A1(_02137_),
    .A2(_07720_),
    .B1(_07731_),
    .B2(_07737_),
    .C1(_08112_),
    .X(_08488_));
 sky130_fd_sc_hd__a21oi_1 _18888_ (.A1(net299),
    .A2(_08106_),
    .B1(_08114_),
    .Y(_08489_));
 sky130_fd_sc_hd__a22oi_2 _18889_ (.A1(_08104_),
    .A2(_08108_),
    .B1(_08114_),
    .B2(_08112_),
    .Y(_08490_));
 sky130_fd_sc_hd__o2bb2ai_1 _18890_ (.A1_N(_08104_),
    .A2_N(_08108_),
    .B1(_08115_),
    .B2(_08111_),
    .Y(_08492_));
 sky130_fd_sc_hd__a31oi_2 _18891_ (.A1(_08482_),
    .A2(_08483_),
    .A3(net312),
    .B1(net293),
    .Y(_08493_));
 sky130_fd_sc_hd__a31o_1 _18892_ (.A1(_08482_),
    .A2(_08483_),
    .A3(net312),
    .B1(net293),
    .X(_08494_));
 sky130_fd_sc_hd__a311oi_4 _18893_ (.A1(_08482_),
    .A2(_08483_),
    .A3(net312),
    .B1(net293),
    .C1(_08472_),
    .Y(_08495_));
 sky130_fd_sc_hd__a2bb2oi_4 _18894_ (.A1_N(_05242_),
    .A2_N(net314),
    .B1(_08473_),
    .B2(_08485_),
    .Y(_08496_));
 sky130_fd_sc_hd__o21ai_1 _18895_ (.A1(_05242_),
    .A2(net314),
    .B1(_08487_),
    .Y(_08497_));
 sky130_fd_sc_hd__o211ai_1 _18896_ (.A1(_08494_),
    .A2(_08472_),
    .B1(_08492_),
    .C1(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__o22ai_1 _18897_ (.A1(_08111_),
    .A2(_08489_),
    .B1(_08495_),
    .B2(_08496_),
    .Y(_08499_));
 sky130_fd_sc_hd__nand3_1 _18898_ (.A(_08498_),
    .B(_08499_),
    .C(net308),
    .Y(_08500_));
 sky130_fd_sc_hd__or3_1 _18899_ (.A(net324),
    .B(_00033_),
    .C(_08486_),
    .X(_08501_));
 sky130_fd_sc_hd__o21ai_1 _18900_ (.A1(net295),
    .A2(_08486_),
    .B1(_08490_),
    .Y(_08503_));
 sky130_fd_sc_hd__o22ai_2 _18901_ (.A1(_08109_),
    .A2(_08488_),
    .B1(_08495_),
    .B2(_08496_),
    .Y(_08504_));
 sky130_fd_sc_hd__o221ai_4 _18902_ (.A1(net324),
    .A2(_00033_),
    .B1(_08495_),
    .B2(_08503_),
    .C1(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__o31a_2 _18903_ (.A1(net324),
    .A2(_00033_),
    .A3(_08486_),
    .B1(_08505_),
    .X(_08506_));
 sky130_fd_sc_hd__o21ai_1 _18904_ (.A1(_01919_),
    .A2(_01930_),
    .B1(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__a2bb2oi_1 _18905_ (.A1_N(_04161_),
    .A2_N(_04184_),
    .B1(_08501_),
    .B2(_08505_),
    .Y(_08508_));
 sky130_fd_sc_hd__o211ai_4 _18906_ (.A1(_08487_),
    .A2(net308),
    .B1(net298),
    .C1(_08500_),
    .Y(_08509_));
 sky130_fd_sc_hd__o211a_1 _18907_ (.A1(net309),
    .A2(_08486_),
    .B1(net299),
    .C1(_08505_),
    .X(_08510_));
 sky130_fd_sc_hd__o211ai_4 _18908_ (.A1(net309),
    .A2(_08486_),
    .B1(net299),
    .C1(_08505_),
    .Y(_08511_));
 sky130_fd_sc_hd__o21ai_2 _18909_ (.A1(_08128_),
    .A2(_08125_),
    .B1(_08124_),
    .Y(_08512_));
 sky130_fd_sc_hd__o2111ai_1 _18910_ (.A1(_08128_),
    .A2(_08125_),
    .B1(_08124_),
    .C1(_08511_),
    .D1(_08509_),
    .Y(_08514_));
 sky130_fd_sc_hd__o22ai_1 _18911_ (.A1(_08123_),
    .A2(_08130_),
    .B1(_08508_),
    .B2(_08510_),
    .Y(_08515_));
 sky130_fd_sc_hd__nand3_1 _18912_ (.A(_08515_),
    .B(net280),
    .C(_08514_),
    .Y(_08516_));
 sky130_fd_sc_hd__o311a_2 _18913_ (.A1(net308),
    .A2(_08472_),
    .A3(_08484_),
    .B1(_08500_),
    .C1(_01973_),
    .X(_08517_));
 sky130_fd_sc_hd__a21oi_4 _18914_ (.A1(_08509_),
    .A2(_08511_),
    .B1(_08512_),
    .Y(_08518_));
 sky130_fd_sc_hd__nand3_2 _18915_ (.A(_08512_),
    .B(_08511_),
    .C(_08509_),
    .Y(_08519_));
 sky130_fd_sc_hd__o21ai_4 _18916_ (.A1(net306),
    .A2(net303),
    .B1(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__o22ai_4 _18917_ (.A1(net280),
    .A2(_08506_),
    .B1(_08518_),
    .B2(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__o22a_2 _18918_ (.A1(net280),
    .A2(_08506_),
    .B1(_08518_),
    .B2(_08520_),
    .X(_08522_));
 sky130_fd_sc_hd__o211ai_4 _18919_ (.A1(_02049_),
    .A2(net342),
    .B1(_08507_),
    .C1(_08516_),
    .Y(_08523_));
 sky130_fd_sc_hd__o22ai_2 _18920_ (.A1(_02093_),
    .A2(_02115_),
    .B1(_08518_),
    .B2(_08520_),
    .Y(_08525_));
 sky130_fd_sc_hd__o221a_1 _18921_ (.A1(net280),
    .A2(_08506_),
    .B1(_08518_),
    .B2(_08520_),
    .C1(_02137_),
    .X(_08526_));
 sky130_fd_sc_hd__o221ai_1 _18922_ (.A1(net280),
    .A2(_08506_),
    .B1(_08518_),
    .B2(_08520_),
    .C1(_02137_),
    .Y(_08527_));
 sky130_fd_sc_hd__o21a_1 _18923_ (.A1(_08517_),
    .A2(_08525_),
    .B1(_08523_),
    .X(_08528_));
 sky130_fd_sc_hd__o21ai_2 _18924_ (.A1(_08517_),
    .A2(_08525_),
    .B1(_08523_),
    .Y(_08529_));
 sky130_fd_sc_hd__and4_1 _18925_ (.A(_07136_),
    .B(_07138_),
    .C(_07422_),
    .D(_07425_),
    .X(_08530_));
 sky130_fd_sc_hd__nand3_1 _18926_ (.A(_07770_),
    .B(_08143_),
    .C(_08530_),
    .Y(_08531_));
 sky130_fd_sc_hd__o211ai_4 _18927_ (.A1(_08147_),
    .A2(_08142_),
    .B1(_08144_),
    .C1(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__nand4_1 _18928_ (.A(_07766_),
    .B(_07769_),
    .C(_08530_),
    .D(_07139_),
    .Y(_08533_));
 sky130_fd_sc_hd__nand3b_4 _18929_ (.A_N(_08533_),
    .B(_08144_),
    .C(_08143_),
    .Y(_08534_));
 sky130_fd_sc_hd__nand2_1 _18930_ (.A(_08532_),
    .B(_08534_),
    .Y(_08536_));
 sky130_fd_sc_hd__a21oi_2 _18931_ (.A1(_08532_),
    .A2(_08534_),
    .B1(_08529_),
    .Y(_08537_));
 sky130_fd_sc_hd__a21o_1 _18932_ (.A1(_08532_),
    .A2(_08534_),
    .B1(_08529_),
    .X(_08538_));
 sky130_fd_sc_hd__a31oi_2 _18933_ (.A1(_08529_),
    .A2(_08532_),
    .A3(_08534_),
    .B1(_04040_),
    .Y(_08539_));
 sky130_fd_sc_hd__o22ai_2 _18934_ (.A1(_04008_),
    .A2(net300),
    .B1(_08528_),
    .B2(_08536_),
    .Y(_08540_));
 sky130_fd_sc_hd__or3_2 _18935_ (.A(_04008_),
    .B(net300),
    .C(_08522_),
    .X(_08541_));
 sky130_fd_sc_hd__inv_2 _18936_ (.A(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__a22o_1 _18937_ (.A1(_08523_),
    .A2(_08527_),
    .B1(_08532_),
    .B2(_08534_),
    .X(_08543_));
 sky130_fd_sc_hd__o211ai_4 _18938_ (.A1(_02148_),
    .A2(_08521_),
    .B1(_08532_),
    .C1(_08534_),
    .Y(_08544_));
 sky130_fd_sc_hd__o2111ai_2 _18939_ (.A1(_02148_),
    .A2(_08521_),
    .B1(_08523_),
    .C1(_08532_),
    .D1(_08534_),
    .Y(_08545_));
 sky130_fd_sc_hd__nand3_2 _18940_ (.A(_08543_),
    .B(_08545_),
    .C(net276),
    .Y(_08547_));
 sky130_fd_sc_hd__a22oi_4 _18941_ (.A1(_04040_),
    .A2(_08522_),
    .B1(_08539_),
    .B2(_08538_),
    .Y(_08548_));
 sky130_fd_sc_hd__inv_2 _18942_ (.A(_08548_),
    .Y(_08549_));
 sky130_fd_sc_hd__o221a_2 _18943_ (.A1(net276),
    .A2(_08521_),
    .B1(_08537_),
    .B2(_08540_),
    .C1(_05234_),
    .X(_08550_));
 sky130_fd_sc_hd__a221o_1 _18944_ (.A1(_04040_),
    .A2(_08522_),
    .B1(_08539_),
    .B2(_08538_),
    .C1(net273),
    .X(_08551_));
 sky130_fd_sc_hd__a31o_1 _18945_ (.A1(_08543_),
    .A2(_08545_),
    .A3(net276),
    .B1(net319),
    .X(_08552_));
 sky130_fd_sc_hd__o311a_1 _18946_ (.A1(_04008_),
    .A2(net300),
    .A3(_08522_),
    .B1(net320),
    .C1(_08547_),
    .X(_08553_));
 sky130_fd_sc_hd__nand3_4 _18947_ (.A(_08547_),
    .B(net320),
    .C(_08541_),
    .Y(_08554_));
 sky130_fd_sc_hd__o221ai_4 _18948_ (.A1(net276),
    .A2(_08521_),
    .B1(_08537_),
    .B2(_08540_),
    .C1(net319),
    .Y(_08555_));
 sky130_fd_sc_hd__o2bb2a_1 _18949_ (.A1_N(net326),
    .A2_N(_08153_),
    .B1(_08155_),
    .B2(_07779_),
    .X(_08556_));
 sky130_fd_sc_hd__o31ai_4 _18950_ (.A1(_07779_),
    .A2(_08155_),
    .A3(_08157_),
    .B1(_08160_),
    .Y(_08558_));
 sky130_fd_sc_hd__o31a_1 _18951_ (.A1(_07779_),
    .A2(_08155_),
    .A3(_08157_),
    .B1(_08160_),
    .X(_08559_));
 sky130_fd_sc_hd__a21oi_1 _18952_ (.A1(_08554_),
    .A2(_08555_),
    .B1(_08558_),
    .Y(_08560_));
 sky130_fd_sc_hd__o2bb2ai_4 _18953_ (.A1_N(_08554_),
    .A2_N(_08555_),
    .B1(_08556_),
    .B2(_08157_),
    .Y(_08561_));
 sky130_fd_sc_hd__nand3_4 _18954_ (.A(_08554_),
    .B(_08555_),
    .C(_08558_),
    .Y(_08562_));
 sky130_fd_sc_hd__a31o_1 _18955_ (.A1(_08554_),
    .A2(_08555_),
    .A3(_08558_),
    .B1(_05234_),
    .X(_08563_));
 sky130_fd_sc_hd__nand3_2 _18956_ (.A(_08561_),
    .B(_08562_),
    .C(net273),
    .Y(_08564_));
 sky130_fd_sc_hd__a31oi_4 _18957_ (.A1(_08561_),
    .A2(_08562_),
    .A3(_05233_),
    .B1(_08550_),
    .Y(_08565_));
 sky130_fd_sc_hd__o22ai_4 _18958_ (.A1(net273),
    .A2(_08549_),
    .B1(_08560_),
    .B2(_08563_),
    .Y(_08566_));
 sky130_fd_sc_hd__a311o_2 _18959_ (.A1(_08561_),
    .A2(_08562_),
    .A3(_05233_),
    .B1(net246),
    .C1(_08550_),
    .X(_08567_));
 sky130_fd_sc_hd__o211a_1 _18960_ (.A1(_07796_),
    .A2(_07798_),
    .B1(_08172_),
    .C1(_07795_),
    .X(_08569_));
 sky130_fd_sc_hd__o221a_1 _18961_ (.A1(net348),
    .A2(_07792_),
    .B1(net330),
    .B2(_08170_),
    .C1(_08177_),
    .X(_08570_));
 sky130_fd_sc_hd__o21ai_2 _18962_ (.A1(_08174_),
    .A2(_08178_),
    .B1(_08172_),
    .Y(_08571_));
 sky130_fd_sc_hd__a311oi_4 _18963_ (.A1(_08561_),
    .A2(_08562_),
    .A3(_05233_),
    .B1(_08550_),
    .C1(net326),
    .Y(_08572_));
 sky130_fd_sc_hd__o221ai_4 _18964_ (.A1(_12867_),
    .A2(_12877_),
    .B1(net273),
    .B2(_08549_),
    .C1(_08564_),
    .Y(_08573_));
 sky130_fd_sc_hd__a2bb2oi_4 _18965_ (.A1_N(_12845_),
    .A2_N(_12856_),
    .B1(_08551_),
    .B2(_08564_),
    .Y(_08574_));
 sky130_fd_sc_hd__o21ai_1 _18966_ (.A1(_12845_),
    .A2(_12856_),
    .B1(_08566_),
    .Y(_08575_));
 sky130_fd_sc_hd__o211ai_2 _18967_ (.A1(_08174_),
    .A2(_08569_),
    .B1(_08573_),
    .C1(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__o22ai_2 _18968_ (.A1(_08171_),
    .A2(_08570_),
    .B1(_08572_),
    .B2(_08574_),
    .Y(_08577_));
 sky130_fd_sc_hd__nand3_4 _18969_ (.A(_08576_),
    .B(_08577_),
    .C(net246),
    .Y(_08578_));
 sky130_fd_sc_hd__or3_1 _18970_ (.A(_05481_),
    .B(net269),
    .C(_08565_),
    .X(_08580_));
 sky130_fd_sc_hd__o21ai_1 _18971_ (.A1(_12888_),
    .A2(_08565_),
    .B1(_08571_),
    .Y(_08581_));
 sky130_fd_sc_hd__o22ai_2 _18972_ (.A1(_08174_),
    .A2(_08569_),
    .B1(_08572_),
    .B2(_08574_),
    .Y(_08582_));
 sky130_fd_sc_hd__o221ai_4 _18973_ (.A1(_05481_),
    .A2(net269),
    .B1(_08572_),
    .B2(_08581_),
    .C1(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__o21ai_2 _18974_ (.A1(net246),
    .A2(_08566_),
    .B1(_08578_),
    .Y(_08584_));
 sky130_fd_sc_hd__and3_2 _18975_ (.A(net330),
    .B(_08567_),
    .C(_08578_),
    .X(_08585_));
 sky130_fd_sc_hd__o211ai_4 _18976_ (.A1(_08566_),
    .A2(net246),
    .B1(net330),
    .C1(_08578_),
    .Y(_08586_));
 sky130_fd_sc_hd__and3_2 _18977_ (.A(_08583_),
    .B(_11298_),
    .C(_08580_),
    .X(_08587_));
 sky130_fd_sc_hd__o211ai_4 _18978_ (.A1(net246),
    .A2(_08565_),
    .B1(_11298_),
    .C1(_08583_),
    .Y(_08588_));
 sky130_fd_sc_hd__a211oi_2 _18979_ (.A1(_07813_),
    .A2(_07815_),
    .B1(_07816_),
    .C1(_08189_),
    .Y(_08589_));
 sky130_fd_sc_hd__o21ai_2 _18980_ (.A1(_08191_),
    .A2(_08194_),
    .B1(_08190_),
    .Y(_08591_));
 sky130_fd_sc_hd__o2bb2ai_4 _18981_ (.A1_N(_08586_),
    .A2_N(_08588_),
    .B1(_08589_),
    .B2(_08191_),
    .Y(_08592_));
 sky130_fd_sc_hd__nand3_2 _18982_ (.A(_08586_),
    .B(_08588_),
    .C(_08591_),
    .Y(_08593_));
 sky130_fd_sc_hd__nand3_2 _18983_ (.A(_08592_),
    .B(_08593_),
    .C(net241),
    .Y(_08594_));
 sky130_fd_sc_hd__and3_2 _18984_ (.A(_05754_),
    .B(_08567_),
    .C(_08578_),
    .X(_08595_));
 sky130_fd_sc_hd__a211o_1 _18985_ (.A1(_08580_),
    .A2(_08583_),
    .B1(net266),
    .C1(_05751_),
    .X(_08596_));
 sky130_fd_sc_hd__a31oi_4 _18986_ (.A1(_08592_),
    .A2(_08593_),
    .A3(net241),
    .B1(_08595_),
    .Y(_08597_));
 sky130_fd_sc_hd__a31o_1 _18987_ (.A1(_08592_),
    .A2(_08593_),
    .A3(net241),
    .B1(_08595_),
    .X(_08598_));
 sky130_fd_sc_hd__a311o_1 _18988_ (.A1(_08592_),
    .A2(_08593_),
    .A3(net241),
    .B1(_08595_),
    .C1(net240),
    .X(_08599_));
 sky130_fd_sc_hd__a22oi_4 _18989_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_08594_),
    .B2(_08596_),
    .Y(_08600_));
 sky130_fd_sc_hd__a22o_1 _18990_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_08594_),
    .B2(_08596_),
    .X(_08602_));
 sky130_fd_sc_hd__o221a_1 _18991_ (.A1(net365),
    .A2(net364),
    .B1(net241),
    .B2(_08584_),
    .C1(_08594_),
    .X(_08603_));
 sky130_fd_sc_hd__a311o_1 _18992_ (.A1(_08592_),
    .A2(_08593_),
    .A3(net241),
    .B1(_08595_),
    .C1(net348),
    .X(_08604_));
 sky130_fd_sc_hd__o21ai_4 _18993_ (.A1(_07828_),
    .A2(_08208_),
    .B1(_08211_),
    .Y(_08605_));
 sky130_fd_sc_hd__o31a_1 _18994_ (.A1(_08863_),
    .A2(_08885_),
    .A3(_08204_),
    .B1(_08605_),
    .X(_08606_));
 sky130_fd_sc_hd__o21ai_4 _18995_ (.A1(_08907_),
    .A2(_08204_),
    .B1(_08605_),
    .Y(_08607_));
 sky130_fd_sc_hd__o21ai_1 _18996_ (.A1(_08600_),
    .A2(_08603_),
    .B1(_08606_),
    .Y(_08608_));
 sky130_fd_sc_hd__a22oi_4 _18997_ (.A1(_08213_),
    .A2(_08605_),
    .B1(_08597_),
    .B2(_10015_),
    .Y(_08609_));
 sky130_fd_sc_hd__a22o_1 _18998_ (.A1(_08213_),
    .A2(_08605_),
    .B1(_08597_),
    .B2(_10015_),
    .X(_08610_));
 sky130_fd_sc_hd__nand3_1 _18999_ (.A(_08602_),
    .B(_08606_),
    .C(_08604_),
    .Y(_08611_));
 sky130_fd_sc_hd__o21ai_1 _19000_ (.A1(_08600_),
    .A2(_08603_),
    .B1(_08607_),
    .Y(_08613_));
 sky130_fd_sc_hd__o211ai_4 _19001_ (.A1(net259),
    .A2(net256),
    .B1(_08611_),
    .C1(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__or3_2 _19002_ (.A(net259),
    .B(net256),
    .C(_08597_),
    .X(_08615_));
 sky130_fd_sc_hd__o221ai_4 _19003_ (.A1(net259),
    .A2(net256),
    .B1(_08600_),
    .B2(_08610_),
    .C1(_08608_),
    .Y(_08616_));
 sky130_fd_sc_hd__o311a_2 _19004_ (.A1(net259),
    .A2(_08598_),
    .A3(net256),
    .B1(_06294_),
    .C1(_08614_),
    .X(_08617_));
 sky130_fd_sc_hd__a22o_1 _19005_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_08615_),
    .B2(_08616_),
    .X(_08618_));
 sky130_fd_sc_hd__nand3_4 _19006_ (.A(_08616_),
    .B(_08907_),
    .C(_08615_),
    .Y(_08619_));
 sky130_fd_sc_hd__o311a_1 _19007_ (.A1(net259),
    .A2(_08598_),
    .A3(net256),
    .B1(_08918_),
    .C1(_08614_),
    .X(_08620_));
 sky130_fd_sc_hd__o211ai_4 _19008_ (.A1(_08819_),
    .A2(_08841_),
    .B1(_08599_),
    .C1(_08614_),
    .Y(_08621_));
 sky130_fd_sc_hd__o21a_1 _19009_ (.A1(_07888_),
    .A2(_08219_),
    .B1(_08221_),
    .X(_08622_));
 sky130_fd_sc_hd__o21ai_1 _19010_ (.A1(_08221_),
    .A2(_08222_),
    .B1(_08225_),
    .Y(_08624_));
 sky130_fd_sc_hd__o2bb2ai_4 _19011_ (.A1_N(_08619_),
    .A2_N(_08621_),
    .B1(_08622_),
    .B2(_08222_),
    .Y(_08625_));
 sky130_fd_sc_hd__o211ai_4 _19012_ (.A1(_08224_),
    .A2(_08231_),
    .B1(_08619_),
    .C1(_08621_),
    .Y(_08626_));
 sky130_fd_sc_hd__nand3_1 _19013_ (.A(_08625_),
    .B(_08626_),
    .C(net212),
    .Y(_08627_));
 sky130_fd_sc_hd__a31oi_2 _19014_ (.A1(_08625_),
    .A2(_08626_),
    .A3(net212),
    .B1(_08617_),
    .Y(_08628_));
 sky130_fd_sc_hd__a31o_2 _19015_ (.A1(_08625_),
    .A2(_08626_),
    .A3(net212),
    .B1(_08617_),
    .X(_08629_));
 sky130_fd_sc_hd__or3_1 _19016_ (.A(_06608_),
    .B(net237),
    .C(_08628_),
    .X(_08630_));
 sky130_fd_sc_hd__a2bb2oi_1 _19017_ (.A1_N(_07800_),
    .A2_N(_07822_),
    .B1(_08618_),
    .B2(_08627_),
    .Y(_08631_));
 sky130_fd_sc_hd__a22o_1 _19018_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_08618_),
    .B2(_08627_),
    .X(_08632_));
 sky130_fd_sc_hd__a311oi_4 _19019_ (.A1(_08625_),
    .A2(_08626_),
    .A3(net212),
    .B1(_08617_),
    .C1(_07899_),
    .Y(_08633_));
 sky130_fd_sc_hd__a311o_1 _19020_ (.A1(_08625_),
    .A2(_08626_),
    .A3(net212),
    .B1(_08617_),
    .C1(_07899_),
    .X(_08635_));
 sky130_fd_sc_hd__a32oi_1 _19021_ (.A1(_08234_),
    .A2(_07033_),
    .A3(_08230_),
    .B1(_07861_),
    .B2(_07869_),
    .Y(_08636_));
 sky130_fd_sc_hd__a21oi_2 _19022_ (.A1(_07925_),
    .A2(_08236_),
    .B1(_08237_),
    .Y(_08637_));
 sky130_fd_sc_hd__o21bai_1 _19023_ (.A1(_08631_),
    .A2(_08633_),
    .B1_N(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__nand3_1 _19024_ (.A(_08632_),
    .B(_08635_),
    .C(_08637_),
    .Y(_08639_));
 sky130_fd_sc_hd__o21ai_1 _19025_ (.A1(_08631_),
    .A2(_08633_),
    .B1(_08637_),
    .Y(_08640_));
 sky130_fd_sc_hd__o221ai_1 _19026_ (.A1(_07899_),
    .A2(_08629_),
    .B1(_08636_),
    .B2(_08237_),
    .C1(_08632_),
    .Y(_08641_));
 sky130_fd_sc_hd__nand3_1 _19027_ (.A(_08640_),
    .B(_08641_),
    .C(net211),
    .Y(_08642_));
 sky130_fd_sc_hd__nand3_2 _19028_ (.A(_08638_),
    .B(_08639_),
    .C(net211),
    .Y(_08643_));
 sky130_fd_sc_hd__o21ai_2 _19029_ (.A1(net211),
    .A2(_08629_),
    .B1(_08643_),
    .Y(_08644_));
 sky130_fd_sc_hd__o311a_1 _19030_ (.A1(_06608_),
    .A2(_08629_),
    .A3(net237),
    .B1(_06904_),
    .C1(_08643_),
    .X(_08646_));
 sky130_fd_sc_hd__or3_1 _19031_ (.A(net230),
    .B(_06901_),
    .C(_08644_),
    .X(_08647_));
 sky130_fd_sc_hd__a21oi_2 _19032_ (.A1(_08249_),
    .A2(_08251_),
    .B1(_08247_),
    .Y(_08648_));
 sky130_fd_sc_hd__a21o_1 _19033_ (.A1(_08249_),
    .A2(_08251_),
    .B1(_08247_),
    .X(_08649_));
 sky130_fd_sc_hd__nand3_4 _19034_ (.A(_08642_),
    .B(_07033_),
    .C(_08630_),
    .Y(_08650_));
 sky130_fd_sc_hd__o211ai_4 _19035_ (.A1(_08629_),
    .A2(net211),
    .B1(_07044_),
    .C1(_08643_),
    .Y(_08651_));
 sky130_fd_sc_hd__nand2_1 _19036_ (.A(_08650_),
    .B(_08651_),
    .Y(_08652_));
 sky130_fd_sc_hd__o211a_1 _19037_ (.A1(_08247_),
    .A2(_08256_),
    .B1(_08650_),
    .C1(_08651_),
    .X(_08653_));
 sky130_fd_sc_hd__o211ai_4 _19038_ (.A1(_08247_),
    .A2(_08256_),
    .B1(_08650_),
    .C1(_08651_),
    .Y(_08654_));
 sky130_fd_sc_hd__a21o_1 _19039_ (.A1(_08650_),
    .A2(_08651_),
    .B1(_08649_),
    .X(_08655_));
 sky130_fd_sc_hd__a221oi_1 _19040_ (.A1(_06900_),
    .A2(_06902_),
    .B1(_08652_),
    .B2(_08648_),
    .C1(_08653_),
    .Y(_08657_));
 sky130_fd_sc_hd__o211ai_2 _19041_ (.A1(net230),
    .A2(_06901_),
    .B1(_08654_),
    .C1(_08655_),
    .Y(_08658_));
 sky130_fd_sc_hd__a211o_2 _19042_ (.A1(_08647_),
    .A2(_08658_),
    .B1(_07227_),
    .C1(net203),
    .X(_08659_));
 sky130_fd_sc_hd__a311oi_4 _19043_ (.A1(_08655_),
    .A2(net208),
    .A3(_08654_),
    .B1(_08646_),
    .C1(_06343_),
    .Y(_08660_));
 sky130_fd_sc_hd__a311o_1 _19044_ (.A1(_08655_),
    .A2(net208),
    .A3(_08654_),
    .B1(_08646_),
    .C1(_06343_),
    .X(_08661_));
 sky130_fd_sc_hd__a2bb2oi_2 _19045_ (.A1_N(net394),
    .A2_N(_06267_),
    .B1(_08647_),
    .B2(_08658_),
    .Y(_08662_));
 sky130_fd_sc_hd__o22ai_1 _19046_ (.A1(net394),
    .A2(_06267_),
    .B1(_08646_),
    .B2(_08657_),
    .Y(_08663_));
 sky130_fd_sc_hd__a31oi_1 _19047_ (.A1(_08246_),
    .A2(_08259_),
    .A3(_08265_),
    .B1(_08264_),
    .Y(_08664_));
 sky130_fd_sc_hd__a31o_1 _19048_ (.A1(_08246_),
    .A2(_08259_),
    .A3(_08265_),
    .B1(_08264_),
    .X(_08665_));
 sky130_fd_sc_hd__nand3_1 _19049_ (.A(_08661_),
    .B(_08663_),
    .C(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__o21ai_1 _19050_ (.A1(_08660_),
    .A2(_08662_),
    .B1(_08664_),
    .Y(_08668_));
 sky130_fd_sc_hd__o211ai_4 _19051_ (.A1(_07227_),
    .A2(net203),
    .B1(_08666_),
    .C1(_08668_),
    .Y(_08669_));
 sky130_fd_sc_hd__o21ai_2 _19052_ (.A1(_08274_),
    .A2(_08270_),
    .B1(_08273_),
    .Y(_08670_));
 sky130_fd_sc_hd__o211a_1 _19053_ (.A1(_08274_),
    .A2(_08270_),
    .B1(_05851_),
    .C1(_08273_),
    .X(_08671_));
 sky130_fd_sc_hd__o21ai_1 _19054_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_08670_),
    .Y(_08672_));
 sky130_fd_sc_hd__a21oi_1 _19055_ (.A1(_05862_),
    .A2(_08670_),
    .B1(_07550_),
    .Y(_08673_));
 sky130_fd_sc_hd__a22o_1 _19056_ (.A1(_07545_),
    .A2(_07547_),
    .B1(_08670_),
    .B2(_05862_),
    .X(_08674_));
 sky130_fd_sc_hd__o2111ai_4 _19057_ (.A1(_05862_),
    .A2(_08670_),
    .B1(_08673_),
    .C1(_08659_),
    .D1(_08669_),
    .Y(_08675_));
 sky130_fd_sc_hd__o2bb2ai_2 _19058_ (.A1_N(_08659_),
    .A2_N(_08669_),
    .B1(_08671_),
    .B2(_08674_),
    .Y(_08676_));
 sky130_fd_sc_hd__nand2_1 _19059_ (.A(_08675_),
    .B(_08676_),
    .Y(_08677_));
 sky130_fd_sc_hd__a32oi_4 _19060_ (.A1(_05250_),
    .A2(_08278_),
    .A3(_08279_),
    .B1(_08282_),
    .B2(_07919_),
    .Y(_08679_));
 sky130_fd_sc_hd__a32o_1 _19061_ (.A1(_05250_),
    .A2(_08278_),
    .A3(_08279_),
    .B1(_08282_),
    .B2(_07919_),
    .X(_08680_));
 sky130_fd_sc_hd__and3_1 _19062_ (.A(_05556_),
    .B(_08284_),
    .C(_08285_),
    .X(_08681_));
 sky130_fd_sc_hd__o2111ai_4 _19063_ (.A1(_03399_),
    .A2(_05491_),
    .B1(net396),
    .C1(_08284_),
    .D1(_08285_),
    .Y(_08682_));
 sky130_fd_sc_hd__a22o_1 _19064_ (.A1(_05512_),
    .A2(net396),
    .B1(_08284_),
    .B2(_08285_),
    .X(_08683_));
 sky130_fd_sc_hd__o221a_1 _19065_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_05556_),
    .B2(_08679_),
    .C1(_08682_),
    .X(_08684_));
 sky130_fd_sc_hd__o221ai_2 _19066_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_05556_),
    .B2(_08679_),
    .C1(_08682_),
    .Y(_08685_));
 sky130_fd_sc_hd__nor2_1 _19067_ (.A(_08677_),
    .B(_08684_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand3_1 _19068_ (.A(_08675_),
    .B(_08676_),
    .C(_08685_),
    .Y(_08687_));
 sky130_fd_sc_hd__and4_1 _19069_ (.A(_08677_),
    .B(_08682_),
    .C(_08683_),
    .D(net160),
    .X(_08688_));
 sky130_fd_sc_hd__nand4_1 _19070_ (.A(_08677_),
    .B(_08682_),
    .C(_08683_),
    .D(net160),
    .Y(_08690_));
 sky130_fd_sc_hd__nand3_1 _19071_ (.A(_08684_),
    .B(_08676_),
    .C(_08675_),
    .Y(_08691_));
 sky130_fd_sc_hd__nand2_1 _19072_ (.A(_08677_),
    .B(_08685_),
    .Y(_08692_));
 sky130_fd_sc_hd__a41o_1 _19073_ (.A1(net160),
    .A2(_08677_),
    .A3(_08682_),
    .A4(_08683_),
    .B1(_08686_),
    .X(_08693_));
 sky130_fd_sc_hd__and3_1 _19074_ (.A(_08687_),
    .B(_08690_),
    .C(_05239_),
    .X(_08694_));
 sky130_fd_sc_hd__a21o_1 _19075_ (.A1(_08691_),
    .A2(_08692_),
    .B1(_05250_),
    .X(_08695_));
 sky130_fd_sc_hd__a21oi_2 _19076_ (.A1(_08687_),
    .A2(_08690_),
    .B1(_05239_),
    .Y(_08696_));
 sky130_fd_sc_hd__o21ai_1 _19077_ (.A1(_08694_),
    .A2(_08696_),
    .B1(_08290_),
    .Y(_08697_));
 sky130_fd_sc_hd__a31oi_2 _19078_ (.A1(_05250_),
    .A2(_08691_),
    .A3(_08692_),
    .B1(_08290_),
    .Y(_08698_));
 sky130_fd_sc_hd__a21oi_1 _19079_ (.A1(_08698_),
    .A2(_08695_),
    .B1(_08301_),
    .Y(_08699_));
 sky130_fd_sc_hd__a2bb2o_1 _19080_ (.A1_N(_08300_),
    .A2_N(_08693_),
    .B1(_08697_),
    .B2(_08699_),
    .X(_08701_));
 sky130_fd_sc_hd__nand2_2 _19081_ (.A(net1),
    .B(_08701_),
    .Y(_08702_));
 sky130_fd_sc_hd__or2_1 _19082_ (.A(net1),
    .B(_08701_),
    .X(_08703_));
 sky130_fd_sc_hd__or2_4 _19083_ (.A(net48),
    .B(_08292_),
    .X(_08704_));
 sky130_fd_sc_hd__and3_4 _19084_ (.A(_08704_),
    .B(net49),
    .C(net409),
    .X(_08705_));
 sky130_fd_sc_hd__o211ai_4 _19085_ (.A1(net48),
    .A2(_08292_),
    .B1(net49),
    .C1(net409),
    .Y(_08706_));
 sky130_fd_sc_hd__a21oi_4 _19086_ (.A1(_08704_),
    .A2(net409),
    .B1(net49),
    .Y(_08707_));
 sky130_fd_sc_hd__a21o_4 _19087_ (.A1(_08704_),
    .A2(net409),
    .B1(net49),
    .X(_08708_));
 sky130_fd_sc_hd__a21boi_4 _19088_ (.A1(_08704_),
    .A2(net409),
    .B1_N(net49),
    .Y(_08709_));
 sky130_fd_sc_hd__a21bo_4 _19089_ (.A1(_08704_),
    .A2(net409),
    .B1_N(net49),
    .X(_08710_));
 sky130_fd_sc_hd__and3b_4 _19090_ (.A_N(net49),
    .B(_08704_),
    .C(net409),
    .X(_08712_));
 sky130_fd_sc_hd__nand3b_4 _19091_ (.A_N(net49),
    .B(_08704_),
    .C(net409),
    .Y(_08713_));
 sky130_fd_sc_hd__nand2_8 _19092_ (.A(_08710_),
    .B(_08713_),
    .Y(_08714_));
 sky130_fd_sc_hd__nand2_8 _19093_ (.A(_08706_),
    .B(_08708_),
    .Y(_08715_));
 sky130_fd_sc_hd__a22o_1 _19094_ (.A1(_08702_),
    .A2(_08703_),
    .B1(_08710_),
    .B2(_08713_),
    .X(_08716_));
 sky130_fd_sc_hd__o21ai_1 _19095_ (.A1(_08701_),
    .A2(_08714_),
    .B1(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__o21ai_1 _19096_ (.A1(_05051_),
    .A2(_08305_),
    .B1(_08717_),
    .Y(_08718_));
 sky130_fd_sc_hd__or3_1 _19097_ (.A(_05051_),
    .B(_08305_),
    .C(_08717_),
    .X(_08719_));
 sky130_fd_sc_hd__and2_1 _19098_ (.A(_08718_),
    .B(_08719_),
    .X(net81));
 sky130_fd_sc_hd__o2bb2a_1 _19099_ (.A1_N(_08305_),
    .A2_N(_08717_),
    .B1(_04832_),
    .B2(_04942_),
    .X(_08720_));
 sky130_fd_sc_hd__o32ai_4 _19100_ (.A1(_07844_),
    .A2(_07866_),
    .A3(_08628_),
    .B1(_08633_),
    .B2(_08637_),
    .Y(_08722_));
 sky130_fd_sc_hd__or4_4 _19101_ (.A(net15),
    .B(net16),
    .C(net17),
    .D(_07554_),
    .X(_08723_));
 sky130_fd_sc_hd__and3b_4 _19102_ (.A_N(net18),
    .B(_08723_),
    .C(net410),
    .X(_08724_));
 sky130_fd_sc_hd__inv_2 _19103_ (.A(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__a21boi_4 _19104_ (.A1(_08723_),
    .A2(net410),
    .B1_N(net18),
    .Y(_08726_));
 sky130_fd_sc_hd__inv_2 _19105_ (.A(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__o311a_4 _19106_ (.A1(net16),
    .A2(net17),
    .A3(_07926_),
    .B1(net18),
    .C1(net410),
    .X(_08728_));
 sky130_fd_sc_hd__a21oi_4 _19107_ (.A1(_08723_),
    .A2(net410),
    .B1(net18),
    .Y(_08729_));
 sky130_fd_sc_hd__nor2_4 _19108_ (.A(_08724_),
    .B(net196),
    .Y(_08730_));
 sky130_fd_sc_hd__nor2_8 _19109_ (.A(_08728_),
    .B(_08729_),
    .Y(_08731_));
 sky130_fd_sc_hd__or3_4 _19110_ (.A(_03178_),
    .B(_08728_),
    .C(net195),
    .X(_08733_));
 sky130_fd_sc_hd__o221a_2 _19111_ (.A1(_05130_),
    .A2(_05152_),
    .B1(_08724_),
    .B2(_08726_),
    .C1(net33),
    .X(_08734_));
 sky130_fd_sc_hd__or4_4 _19112_ (.A(_07253_),
    .B(_07572_),
    .C(_07943_),
    .D(_08320_),
    .X(_08735_));
 sky130_fd_sc_hd__inv_2 _19113_ (.A(_08735_),
    .Y(_08736_));
 sky130_fd_sc_hd__o31a_1 _19114_ (.A1(_03178_),
    .A2(_07935_),
    .A3(net199),
    .B1(_08735_),
    .X(_08737_));
 sky130_fd_sc_hd__nand2_1 _19115_ (.A(_08324_),
    .B(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__a22oi_4 _19116_ (.A1(_07254_),
    .A2(_08736_),
    .B1(_08324_),
    .B2(_08737_),
    .Y(_08739_));
 sky130_fd_sc_hd__o2bb2ai_1 _19117_ (.A1_N(_08737_),
    .A2_N(_08324_),
    .B1(_07255_),
    .B2(_08735_),
    .Y(_08740_));
 sky130_fd_sc_hd__a211o_1 _19118_ (.A1(net175),
    .A2(net33),
    .B1(_08307_),
    .C1(_08309_),
    .X(_08741_));
 sky130_fd_sc_hd__or4_1 _19119_ (.A(_03178_),
    .B(_08311_),
    .C(_08312_),
    .D(net177),
    .X(_08742_));
 sky130_fd_sc_hd__o31a_2 _19120_ (.A1(_08728_),
    .A2(net195),
    .A3(_08317_),
    .B1(_08741_),
    .X(_08744_));
 sky130_fd_sc_hd__o21ai_2 _19121_ (.A1(_08317_),
    .A2(net177),
    .B1(_08741_),
    .Y(_08745_));
 sky130_fd_sc_hd__nand2_2 _19122_ (.A(_08740_),
    .B(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__o211ai_4 _19123_ (.A1(_07255_),
    .A2(_08735_),
    .B1(_08744_),
    .C1(_08738_),
    .Y(_08747_));
 sky130_fd_sc_hd__a31oi_4 _19124_ (.A1(_08746_),
    .A2(_08747_),
    .A3(net405),
    .B1(_08734_),
    .Y(_08748_));
 sky130_fd_sc_hd__or3_1 _19125_ (.A(_05348_),
    .B(net401),
    .C(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__a311oi_4 _19126_ (.A1(_08746_),
    .A2(_08747_),
    .A3(net405),
    .B1(_07936_),
    .C1(_08734_),
    .Y(_08750_));
 sky130_fd_sc_hd__a311o_1 _19127_ (.A1(_08746_),
    .A2(_08747_),
    .A3(net405),
    .B1(_07936_),
    .C1(_08734_),
    .X(_08751_));
 sky130_fd_sc_hd__a21oi_2 _19128_ (.A1(_07929_),
    .A2(_07932_),
    .B1(_08748_),
    .Y(_08752_));
 sky130_fd_sc_hd__a21o_1 _19129_ (.A1(_07929_),
    .A2(_07932_),
    .B1(_08748_),
    .X(_08753_));
 sky130_fd_sc_hd__nor2_1 _19130_ (.A(_08750_),
    .B(_08752_),
    .Y(_08755_));
 sky130_fd_sc_hd__nand2_1 _19131_ (.A(_08751_),
    .B(_08753_),
    .Y(_08756_));
 sky130_fd_sc_hd__a22oi_1 _19132_ (.A1(_08327_),
    .A2(_08331_),
    .B1(_08336_),
    .B2(_08330_),
    .Y(_08757_));
 sky130_fd_sc_hd__o22ai_2 _19133_ (.A1(_08325_),
    .A2(_08332_),
    .B1(_08334_),
    .B2(_08335_),
    .Y(_08758_));
 sky130_fd_sc_hd__nand2_1 _19134_ (.A(_08758_),
    .B(_08755_),
    .Y(_08759_));
 sky130_fd_sc_hd__o221ai_4 _19135_ (.A1(_08750_),
    .A2(_08752_),
    .B1(_08334_),
    .B2(_08335_),
    .C1(_08333_),
    .Y(_08760_));
 sky130_fd_sc_hd__o211ai_4 _19136_ (.A1(_05348_),
    .A2(net401),
    .B1(_08759_),
    .C1(_08760_),
    .Y(_08761_));
 sky130_fd_sc_hd__and3_1 _19137_ (.A(_08748_),
    .B(_05381_),
    .C(_05359_),
    .X(_08762_));
 sky130_fd_sc_hd__a21oi_2 _19138_ (.A1(_08759_),
    .A2(_08760_),
    .B1(_05392_),
    .Y(_08763_));
 sky130_fd_sc_hd__o21a_1 _19139_ (.A1(_05403_),
    .A2(_08748_),
    .B1(_08761_),
    .X(_08764_));
 sky130_fd_sc_hd__or4_2 _19140_ (.A(_05676_),
    .B(_05698_),
    .C(_08762_),
    .D(_08763_),
    .X(_08766_));
 sky130_fd_sc_hd__a2bb2oi_1 _19141_ (.A1_N(_07555_),
    .A2_N(net218),
    .B1(_08749_),
    .B2(_08761_),
    .Y(_08767_));
 sky130_fd_sc_hd__a22o_2 _19142_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_08749_),
    .B2(_08761_),
    .X(_08768_));
 sky130_fd_sc_hd__o211ai_4 _19143_ (.A1(_05403_),
    .A2(_08748_),
    .B1(_07564_),
    .C1(_08761_),
    .Y(_08769_));
 sky130_fd_sc_hd__o41a_1 _19144_ (.A1(_07560_),
    .A2(_07562_),
    .A3(_08762_),
    .A4(_08763_),
    .B1(_08769_),
    .X(_08770_));
 sky130_fd_sc_hd__nand2_4 _19145_ (.A(_08768_),
    .B(_08769_),
    .Y(_08771_));
 sky130_fd_sc_hd__a21oi_4 _19146_ (.A1(_08355_),
    .A2(_08352_),
    .B1(_08349_),
    .Y(_08772_));
 sky130_fd_sc_hd__o32ai_1 _19147_ (.A1(net224),
    .A2(_08343_),
    .A3(_08344_),
    .B1(_08353_),
    .B2(_08354_),
    .Y(_08773_));
 sky130_fd_sc_hd__o21ai_1 _19148_ (.A1(_08349_),
    .A2(_08356_),
    .B1(_08770_),
    .Y(_08774_));
 sky130_fd_sc_hd__o311a_2 _19149_ (.A1(net224),
    .A2(_08343_),
    .A3(_08344_),
    .B1(_08357_),
    .C1(_08771_),
    .X(_08775_));
 sky130_fd_sc_hd__o211ai_1 _19150_ (.A1(net224),
    .A2(_08345_),
    .B1(_08357_),
    .C1(_08771_),
    .Y(_08777_));
 sky130_fd_sc_hd__o22ai_4 _19151_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_08771_),
    .B2(_08772_),
    .Y(_08778_));
 sky130_fd_sc_hd__nand3_1 _19152_ (.A(_08774_),
    .B(_08777_),
    .C(net358),
    .Y(_08779_));
 sky130_fd_sc_hd__o22a_1 _19153_ (.A1(net358),
    .A2(_08764_),
    .B1(_08775_),
    .B2(_08778_),
    .X(_08780_));
 sky130_fd_sc_hd__o22ai_2 _19154_ (.A1(net358),
    .A2(_08764_),
    .B1(_08775_),
    .B2(_08778_),
    .Y(_08781_));
 sky130_fd_sc_hd__and3_1 _19155_ (.A(_06804_),
    .B(_06826_),
    .C(_08781_),
    .X(_08782_));
 sky130_fd_sc_hd__or3_2 _19156_ (.A(_06793_),
    .B(_06815_),
    .C(_08780_),
    .X(_08783_));
 sky130_fd_sc_hd__a2bb2oi_2 _19157_ (.A1_N(_07242_),
    .A2_N(_07243_),
    .B1(_08766_),
    .B2(_08779_),
    .Y(_08784_));
 sky130_fd_sc_hd__o21ai_4 _19158_ (.A1(_07242_),
    .A2(_07243_),
    .B1(_08781_),
    .Y(_08785_));
 sky130_fd_sc_hd__o22a_1 _19159_ (.A1(_07244_),
    .A2(_07245_),
    .B1(_08775_),
    .B2(_08778_),
    .X(_08786_));
 sky130_fd_sc_hd__o221ai_4 _19160_ (.A1(net358),
    .A2(_08764_),
    .B1(_08775_),
    .B2(_08778_),
    .C1(net224),
    .Y(_08787_));
 sky130_fd_sc_hd__a21oi_4 _19161_ (.A1(_08766_),
    .A2(_08786_),
    .B1(_08784_),
    .Y(_08788_));
 sky130_fd_sc_hd__nand2_4 _19162_ (.A(_08785_),
    .B(_08787_),
    .Y(_08789_));
 sky130_fd_sc_hd__a31oi_4 _19163_ (.A1(_08371_),
    .A2(_08377_),
    .A3(_08380_),
    .B1(_08365_),
    .Y(_08790_));
 sky130_fd_sc_hd__o22ai_4 _19164_ (.A1(net227),
    .A2(_08362_),
    .B1(_08384_),
    .B2(_08376_),
    .Y(_08791_));
 sky130_fd_sc_hd__a21oi_1 _19165_ (.A1(_08366_),
    .A2(_08385_),
    .B1(_08789_),
    .Y(_08792_));
 sky130_fd_sc_hd__nand2_2 _19166_ (.A(_08791_),
    .B(_08788_),
    .Y(_08793_));
 sky130_fd_sc_hd__o211ai_2 _19167_ (.A1(net227),
    .A2(_08362_),
    .B1(_08385_),
    .C1(_08789_),
    .Y(_08794_));
 sky130_fd_sc_hd__o22ai_1 _19168_ (.A1(net379),
    .A2(net378),
    .B1(_08788_),
    .B2(_08791_),
    .Y(_08795_));
 sky130_fd_sc_hd__o221ai_4 _19169_ (.A1(net379),
    .A2(net378),
    .B1(_08788_),
    .B2(_08791_),
    .C1(_08793_),
    .Y(_08796_));
 sky130_fd_sc_hd__o22a_1 _19170_ (.A1(net357),
    .A2(_08780_),
    .B1(_08792_),
    .B2(_08795_),
    .X(_08798_));
 sky130_fd_sc_hd__a31o_2 _19171_ (.A1(_08793_),
    .A2(_08794_),
    .A3(net357),
    .B1(_08782_),
    .X(_08799_));
 sky130_fd_sc_hd__a2bb2oi_2 _19172_ (.A1_N(_06914_),
    .A2_N(_06916_),
    .B1(_08783_),
    .B2(_08796_),
    .Y(_08800_));
 sky130_fd_sc_hd__a22o_1 _19173_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_08783_),
    .B2(_08796_),
    .X(_08801_));
 sky130_fd_sc_hd__a31oi_1 _19174_ (.A1(_08793_),
    .A2(_08794_),
    .A3(net357),
    .B1(net225),
    .Y(_08802_));
 sky130_fd_sc_hd__o221a_2 _19175_ (.A1(net357),
    .A2(_08780_),
    .B1(_08792_),
    .B2(_08795_),
    .C1(net227),
    .X(_08803_));
 sky130_fd_sc_hd__a311o_1 _19176_ (.A1(_08793_),
    .A2(_08794_),
    .A3(net357),
    .B1(net225),
    .C1(_08782_),
    .X(_08804_));
 sky130_fd_sc_hd__a21oi_2 _19177_ (.A1(_08783_),
    .A2(_08802_),
    .B1(_08800_),
    .Y(_08805_));
 sky130_fd_sc_hd__and3_1 _19178_ (.A(_07637_),
    .B(_07639_),
    .C(_07311_),
    .X(_08806_));
 sky130_fd_sc_hd__nand4_1 _19179_ (.A(_08806_),
    .B(_08012_),
    .C(_08009_),
    .D(_07313_),
    .Y(_08807_));
 sky130_fd_sc_hd__nand3_1 _19180_ (.A(_08399_),
    .B(_08806_),
    .C(_08013_),
    .Y(_08809_));
 sky130_fd_sc_hd__nor3_2 _19181_ (.A(_08807_),
    .B(_08400_),
    .C(_08398_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand3b_2 _19182_ (.A_N(_08807_),
    .B(_08401_),
    .C(_08399_),
    .Y(_08811_));
 sky130_fd_sc_hd__o211a_1 _19183_ (.A1(_08396_),
    .A2(_08398_),
    .B1(_08401_),
    .C1(_08809_),
    .X(_08812_));
 sky130_fd_sc_hd__o211ai_4 _19184_ (.A1(_08396_),
    .A2(_08398_),
    .B1(_08401_),
    .C1(_08809_),
    .Y(_08813_));
 sky130_fd_sc_hd__nand2_2 _19185_ (.A(_08811_),
    .B(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__o21ai_1 _19186_ (.A1(_08810_),
    .A2(_08812_),
    .B1(_08805_),
    .Y(_08815_));
 sky130_fd_sc_hd__nand4_4 _19187_ (.A(_08801_),
    .B(_08804_),
    .C(_08811_),
    .D(_08813_),
    .Y(_08816_));
 sky130_fd_sc_hd__o22ai_4 _19188_ (.A1(_08800_),
    .A2(_08803_),
    .B1(_08810_),
    .B2(_08812_),
    .Y(_08817_));
 sky130_fd_sc_hd__o221ai_4 _19189_ (.A1(_07691_),
    .A2(net371),
    .B1(_08805_),
    .B2(_08814_),
    .C1(_08815_),
    .Y(_08818_));
 sky130_fd_sc_hd__nand3_2 _19190_ (.A(_08817_),
    .B(net354),
    .C(_08816_),
    .Y(_08820_));
 sky130_fd_sc_hd__a21oi_2 _19191_ (.A1(_08783_),
    .A2(_08796_),
    .B1(net355),
    .Y(_08821_));
 sky130_fd_sc_hd__or3_2 _19192_ (.A(_07691_),
    .B(net371),
    .C(_08798_),
    .X(_08822_));
 sky130_fd_sc_hd__o211a_1 _19193_ (.A1(_08799_),
    .A2(net354),
    .B1(_08732_),
    .C1(_08818_),
    .X(_08823_));
 sky130_fd_sc_hd__a211o_2 _19194_ (.A1(_08820_),
    .A2(_08822_),
    .B1(net353),
    .C1(net352),
    .X(_08824_));
 sky130_fd_sc_hd__a21oi_1 _19195_ (.A1(_08031_),
    .A2(_08419_),
    .B1(_08411_),
    .Y(_08825_));
 sky130_fd_sc_hd__o211a_1 _19196_ (.A1(_08025_),
    .A2(net253),
    .B1(_08419_),
    .C1(_08417_),
    .X(_08826_));
 sky130_fd_sc_hd__a31oi_4 _19197_ (.A1(_08031_),
    .A2(_08417_),
    .A3(_08419_),
    .B1(_08411_),
    .Y(_08827_));
 sky130_fd_sc_hd__a311oi_4 _19198_ (.A1(_08817_),
    .A2(net354),
    .A3(_08816_),
    .B1(_08821_),
    .C1(net232),
    .Y(_08828_));
 sky130_fd_sc_hd__nand3_4 _19199_ (.A(_08820_),
    .B(_08822_),
    .C(net234),
    .Y(_08829_));
 sky130_fd_sc_hd__a21oi_2 _19200_ (.A1(_08820_),
    .A2(_08822_),
    .B1(net234),
    .Y(_08831_));
 sky130_fd_sc_hd__o211ai_4 _19201_ (.A1(_08799_),
    .A2(net354),
    .B1(net232),
    .C1(_08818_),
    .Y(_08832_));
 sky130_fd_sc_hd__o211a_1 _19202_ (.A1(_08411_),
    .A2(_08826_),
    .B1(_08829_),
    .C1(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__o211ai_4 _19203_ (.A1(_08411_),
    .A2(_08826_),
    .B1(_08829_),
    .C1(_08832_),
    .Y(_08834_));
 sky130_fd_sc_hd__a21boi_1 _19204_ (.A1(_08829_),
    .A2(_08832_),
    .B1_N(_08827_),
    .Y(_08835_));
 sky130_fd_sc_hd__o22ai_4 _19205_ (.A1(_08416_),
    .A2(_08825_),
    .B1(_08828_),
    .B2(_08831_),
    .Y(_08836_));
 sky130_fd_sc_hd__nand3_2 _19206_ (.A(_08836_),
    .B(net338),
    .C(_08834_),
    .Y(_08837_));
 sky130_fd_sc_hd__a311o_1 _19207_ (.A1(_08817_),
    .A2(net354),
    .A3(_08816_),
    .B1(_08821_),
    .C1(net338),
    .X(_08838_));
 sky130_fd_sc_hd__o22ai_2 _19208_ (.A1(net353),
    .A2(net352),
    .B1(_08833_),
    .B2(_08835_),
    .Y(_08839_));
 sky130_fd_sc_hd__a31o_1 _19209_ (.A1(_08836_),
    .A2(net338),
    .A3(_08834_),
    .B1(_08823_),
    .X(_08840_));
 sky130_fd_sc_hd__o211ai_4 _19210_ (.A1(_08042_),
    .A2(net262),
    .B1(_08432_),
    .C1(_08060_),
    .Y(_08842_));
 sky130_fd_sc_hd__o211ai_4 _19211_ (.A1(net261),
    .A2(_08043_),
    .B1(_08433_),
    .C1(_08435_),
    .Y(_08843_));
 sky130_fd_sc_hd__a311oi_4 _19212_ (.A1(_08836_),
    .A2(net338),
    .A3(_08834_),
    .B1(net251),
    .C1(_08823_),
    .Y(_08844_));
 sky130_fd_sc_hd__o211ai_4 _19213_ (.A1(_06309_),
    .A2(_06312_),
    .B1(_08824_),
    .C1(_08837_),
    .Y(_08845_));
 sky130_fd_sc_hd__a2bb2oi_4 _19214_ (.A1_N(_06305_),
    .A2_N(net283),
    .B1(_08824_),
    .B2(_08837_),
    .Y(_08846_));
 sky130_fd_sc_hd__o211ai_4 _19215_ (.A1(_06305_),
    .A2(net283),
    .B1(_08838_),
    .C1(_08839_),
    .Y(_08847_));
 sky130_fd_sc_hd__nor2_1 _19216_ (.A(_08844_),
    .B(_08846_),
    .Y(_08848_));
 sky130_fd_sc_hd__o2111ai_4 _19217_ (.A1(_08431_),
    .A2(net254),
    .B1(_08845_),
    .C1(_08843_),
    .D1(_08847_),
    .Y(_08849_));
 sky130_fd_sc_hd__o2bb2ai_1 _19218_ (.A1_N(_08432_),
    .A2_N(_08843_),
    .B1(_08844_),
    .B2(_08846_),
    .Y(_08850_));
 sky130_fd_sc_hd__o211ai_4 _19219_ (.A1(_09785_),
    .A2(_09807_),
    .B1(_08849_),
    .C1(_08850_),
    .Y(_08851_));
 sky130_fd_sc_hd__a211o_1 _19220_ (.A1(_08824_),
    .A2(_08837_),
    .B1(_09785_),
    .C1(_09807_),
    .X(_08853_));
 sky130_fd_sc_hd__o2111ai_1 _19221_ (.A1(net253),
    .A2(_08430_),
    .B1(_08842_),
    .C1(_08845_),
    .D1(_08847_),
    .Y(_08854_));
 sky130_fd_sc_hd__o2bb2ai_1 _19222_ (.A1_N(_08433_),
    .A2_N(_08842_),
    .B1(_08844_),
    .B2(_08846_),
    .Y(_08855_));
 sky130_fd_sc_hd__o211ai_1 _19223_ (.A1(_09785_),
    .A2(_09807_),
    .B1(_08854_),
    .C1(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__o21ai_4 _19224_ (.A1(net336),
    .A2(_08840_),
    .B1(_08851_),
    .Y(_08857_));
 sky130_fd_sc_hd__o211a_1 _19225_ (.A1(_08840_),
    .A2(net336),
    .B1(_11079_),
    .C1(_08851_),
    .X(_08858_));
 sky130_fd_sc_hd__or3_1 _19226_ (.A(_11046_),
    .B(_11057_),
    .C(_08857_),
    .X(_08859_));
 sky130_fd_sc_hd__o211ai_2 _19227_ (.A1(_08840_),
    .A2(net336),
    .B1(net253),
    .C1(_08851_),
    .Y(_08860_));
 sky130_fd_sc_hd__o211ai_2 _19228_ (.A1(net286),
    .A2(_06012_),
    .B1(_08853_),
    .C1(_08856_),
    .Y(_08861_));
 sky130_fd_sc_hd__nand2_4 _19229_ (.A(_08860_),
    .B(_08861_),
    .Y(_08862_));
 sky130_fd_sc_hd__a31oi_4 _19230_ (.A1(_08450_),
    .A2(_08453_),
    .A3(_08461_),
    .B1(_08456_),
    .Y(_08864_));
 sky130_fd_sc_hd__o211ai_2 _19231_ (.A1(net262),
    .A2(_08445_),
    .B1(_08467_),
    .C1(_08862_),
    .Y(_08865_));
 sky130_fd_sc_hd__o211a_1 _19232_ (.A1(_08862_),
    .A2(_08864_),
    .B1(net333),
    .C1(_08865_),
    .X(_08866_));
 sky130_fd_sc_hd__o211ai_4 _19233_ (.A1(_08862_),
    .A2(_08864_),
    .B1(net333),
    .C1(_08865_),
    .Y(_08867_));
 sky130_fd_sc_hd__o21ai_4 _19234_ (.A1(net333),
    .A2(_08857_),
    .B1(_08867_),
    .Y(_08868_));
 sky130_fd_sc_hd__inv_2 _19235_ (.A(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__a2bb2oi_1 _19236_ (.A1_N(_05760_),
    .A2_N(net290),
    .B1(_08859_),
    .B2(_08867_),
    .Y(_08870_));
 sky130_fd_sc_hd__o22ai_2 _19237_ (.A1(_05760_),
    .A2(net290),
    .B1(_08858_),
    .B2(_08866_),
    .Y(_08871_));
 sky130_fd_sc_hd__o211a_1 _19238_ (.A1(net333),
    .A2(_08857_),
    .B1(net262),
    .C1(_08867_),
    .X(_08872_));
 sky130_fd_sc_hd__o211ai_4 _19239_ (.A1(net333),
    .A2(_08857_),
    .B1(net262),
    .C1(_08867_),
    .Y(_08873_));
 sky130_fd_sc_hd__nor2_1 _19240_ (.A(_08870_),
    .B(_08872_),
    .Y(_08875_));
 sky130_fd_sc_hd__nand2_1 _19241_ (.A(_08871_),
    .B(_08873_),
    .Y(_08876_));
 sky130_fd_sc_hd__nand4_2 _19242_ (.A(_07380_),
    .B(_07382_),
    .C(_07709_),
    .D(_07711_),
    .Y(_08877_));
 sky130_fd_sc_hd__a21oi_1 _19243_ (.A1(net293),
    .A2(_08087_),
    .B1(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__a211oi_2 _19244_ (.A1(_08070_),
    .A2(_08091_),
    .B1(_08877_),
    .C1(_08094_),
    .Y(_08879_));
 sky130_fd_sc_hd__o211ai_4 _19245_ (.A1(net293),
    .A2(_08087_),
    .B1(_08878_),
    .C1(_08475_),
    .Y(_08880_));
 sky130_fd_sc_hd__o211a_1 _19246_ (.A1(_08481_),
    .A2(_08474_),
    .B1(_08477_),
    .C1(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__o211ai_4 _19247_ (.A1(_08481_),
    .A2(_08474_),
    .B1(_08477_),
    .C1(_08880_),
    .Y(_08882_));
 sky130_fd_sc_hd__nand4_4 _19248_ (.A(_08879_),
    .B(_08477_),
    .C(_08475_),
    .D(_07378_),
    .Y(_08883_));
 sky130_fd_sc_hd__inv_2 _19249_ (.A(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__o31a_2 _19250_ (.A1(_07377_),
    .A2(_08476_),
    .A3(_08880_),
    .B1(_08882_),
    .X(_08886_));
 sky130_fd_sc_hd__a21oi_2 _19251_ (.A1(_08882_),
    .A2(_08883_),
    .B1(_08876_),
    .Y(_08887_));
 sky130_fd_sc_hd__o211ai_1 _19252_ (.A1(_08870_),
    .A2(_08872_),
    .B1(_08882_),
    .C1(_08883_),
    .Y(_08888_));
 sky130_fd_sc_hd__o21ai_2 _19253_ (.A1(_12670_),
    .A2(net327),
    .B1(_08888_),
    .Y(_08889_));
 sky130_fd_sc_hd__nand4_2 _19254_ (.A(_08871_),
    .B(_08873_),
    .C(_08882_),
    .D(_08883_),
    .Y(_08890_));
 sky130_fd_sc_hd__a22o_1 _19255_ (.A1(_08871_),
    .A2(_08873_),
    .B1(_08882_),
    .B2(_08883_),
    .X(_08891_));
 sky130_fd_sc_hd__a211o_2 _19256_ (.A1(_08859_),
    .A2(_08867_),
    .B1(_12670_),
    .C1(net327),
    .X(_08892_));
 sky130_fd_sc_hd__inv_2 _19257_ (.A(_08892_),
    .Y(_08893_));
 sky130_fd_sc_hd__nand3_1 _19258_ (.A(_08891_),
    .B(net312),
    .C(_08890_),
    .Y(_08894_));
 sky130_fd_sc_hd__a31o_1 _19259_ (.A1(_08891_),
    .A2(net312),
    .A3(_08890_),
    .B1(_08893_),
    .X(_08895_));
 sky130_fd_sc_hd__a311oi_4 _19260_ (.A1(_08891_),
    .A2(net312),
    .A3(_08890_),
    .B1(_08893_),
    .C1(net291),
    .Y(_08897_));
 sky130_fd_sc_hd__nand3_4 _19261_ (.A(_08894_),
    .B(net267),
    .C(_08892_),
    .Y(_08898_));
 sky130_fd_sc_hd__o221ai_4 _19262_ (.A1(net312),
    .A2(_08868_),
    .B1(_08887_),
    .B2(_08889_),
    .C1(net291),
    .Y(_08899_));
 sky130_fd_sc_hd__o221a_1 _19263_ (.A1(_08109_),
    .A2(_08114_),
    .B1(_08486_),
    .B2(net295),
    .C1(_08112_),
    .X(_08900_));
 sky130_fd_sc_hd__o31a_1 _19264_ (.A1(net293),
    .A2(_08472_),
    .A3(_08484_),
    .B1(_08490_),
    .X(_08901_));
 sky130_fd_sc_hd__o32a_1 _19265_ (.A1(_05242_),
    .A2(net314),
    .A3(_08487_),
    .B1(_08490_),
    .B2(_08496_),
    .X(_08902_));
 sky130_fd_sc_hd__o21a_1 _19266_ (.A1(_08495_),
    .A2(_08492_),
    .B1(_08497_),
    .X(_08903_));
 sky130_fd_sc_hd__a21oi_1 _19267_ (.A1(_08898_),
    .A2(_08899_),
    .B1(_08902_),
    .Y(_08904_));
 sky130_fd_sc_hd__o2bb2ai_4 _19268_ (.A1_N(_08898_),
    .A2_N(_08899_),
    .B1(_08900_),
    .B2(_08495_),
    .Y(_08905_));
 sky130_fd_sc_hd__o211a_1 _19269_ (.A1(_08496_),
    .A2(_08901_),
    .B1(_08899_),
    .C1(_08898_),
    .X(_08906_));
 sky130_fd_sc_hd__nand3_4 _19270_ (.A(_08898_),
    .B(_08899_),
    .C(_08902_),
    .Y(_08908_));
 sky130_fd_sc_hd__nand3_2 _19271_ (.A(_08905_),
    .B(_08908_),
    .C(net309),
    .Y(_08909_));
 sky130_fd_sc_hd__o221a_4 _19272_ (.A1(net312),
    .A2(_08868_),
    .B1(_08887_),
    .B2(_08889_),
    .C1(_00066_),
    .X(_08910_));
 sky130_fd_sc_hd__a211o_2 _19273_ (.A1(_08892_),
    .A2(_08894_),
    .B1(net324),
    .C1(_00033_),
    .X(_08911_));
 sky130_fd_sc_hd__o22ai_2 _19274_ (.A1(net324),
    .A2(_00033_),
    .B1(_08904_),
    .B2(_08906_),
    .Y(_08912_));
 sky130_fd_sc_hd__a31oi_4 _19275_ (.A1(_08905_),
    .A2(_08908_),
    .A3(net309),
    .B1(_08910_),
    .Y(_08913_));
 sky130_fd_sc_hd__a31o_1 _19276_ (.A1(_08905_),
    .A2(_08908_),
    .A3(net309),
    .B1(_08910_),
    .X(_08914_));
 sky130_fd_sc_hd__o211a_1 _19277_ (.A1(_08128_),
    .A2(_08125_),
    .B1(_08124_),
    .C1(_08509_),
    .X(_08915_));
 sky130_fd_sc_hd__a21o_1 _19278_ (.A1(_08512_),
    .A2(_08511_),
    .B1(_08508_),
    .X(_08916_));
 sky130_fd_sc_hd__a311oi_4 _19279_ (.A1(_08905_),
    .A2(_08908_),
    .A3(net309),
    .B1(_08910_),
    .C1(net293),
    .Y(_08917_));
 sky130_fd_sc_hd__nand4_2 _19280_ (.A(_05243_),
    .B(_05245_),
    .C(_08909_),
    .D(_08911_),
    .Y(_08919_));
 sky130_fd_sc_hd__a22oi_4 _19281_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_08909_),
    .B2(_08911_),
    .Y(_08920_));
 sky130_fd_sc_hd__o221ai_4 _19282_ (.A1(_05242_),
    .A2(net314),
    .B1(_08895_),
    .B2(net308),
    .C1(_08912_),
    .Y(_08921_));
 sky130_fd_sc_hd__nor2_1 _19283_ (.A(_08917_),
    .B(_08920_),
    .Y(_08922_));
 sky130_fd_sc_hd__o2111ai_1 _19284_ (.A1(net299),
    .A2(_08506_),
    .B1(_08519_),
    .C1(_08919_),
    .D1(_08921_),
    .Y(_08923_));
 sky130_fd_sc_hd__o21ai_1 _19285_ (.A1(_08917_),
    .A2(_08920_),
    .B1(_08916_),
    .Y(_08924_));
 sky130_fd_sc_hd__o211ai_2 _19286_ (.A1(net306),
    .A2(net303),
    .B1(_08923_),
    .C1(_08924_),
    .Y(_08925_));
 sky130_fd_sc_hd__or3_1 _19287_ (.A(net306),
    .B(net303),
    .C(_08913_),
    .X(_08926_));
 sky130_fd_sc_hd__o21ai_1 _19288_ (.A1(net295),
    .A2(_08913_),
    .B1(_08916_),
    .Y(_08927_));
 sky130_fd_sc_hd__o22ai_2 _19289_ (.A1(_08510_),
    .A2(_08915_),
    .B1(_08917_),
    .B2(_08920_),
    .Y(_08928_));
 sky130_fd_sc_hd__o221ai_4 _19290_ (.A1(net306),
    .A2(net303),
    .B1(_08917_),
    .B2(_08927_),
    .C1(_08928_),
    .Y(_08930_));
 sky130_fd_sc_hd__o21ai_2 _19291_ (.A1(net280),
    .A2(_08913_),
    .B1(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__inv_2 _19292_ (.A(_08931_),
    .Y(_08932_));
 sky130_fd_sc_hd__or3_1 _19293_ (.A(_04008_),
    .B(net300),
    .C(_08931_),
    .X(_08933_));
 sky130_fd_sc_hd__a2bb2oi_1 _19294_ (.A1_N(_04161_),
    .A2_N(_04184_),
    .B1(_08926_),
    .B2(_08930_),
    .Y(_08934_));
 sky130_fd_sc_hd__o211ai_4 _19295_ (.A1(_08914_),
    .A2(net280),
    .B1(net298),
    .C1(_08925_),
    .Y(_08935_));
 sky130_fd_sc_hd__o211a_1 _19296_ (.A1(net280),
    .A2(_08913_),
    .B1(net299),
    .C1(_08930_),
    .X(_08936_));
 sky130_fd_sc_hd__o211ai_4 _19297_ (.A1(net280),
    .A2(_08913_),
    .B1(net299),
    .C1(_08930_),
    .Y(_08937_));
 sky130_fd_sc_hd__a22oi_1 _19298_ (.A1(_02148_),
    .A2(_08521_),
    .B1(_08532_),
    .B2(_08534_),
    .Y(_08938_));
 sky130_fd_sc_hd__o2bb2ai_2 _19299_ (.A1_N(_08532_),
    .A2_N(_08534_),
    .B1(_02137_),
    .B2(_08522_),
    .Y(_08939_));
 sky130_fd_sc_hd__o2111ai_1 _19300_ (.A1(_02137_),
    .A2(_08522_),
    .B1(_08544_),
    .C1(_08935_),
    .D1(_08937_),
    .Y(_08941_));
 sky130_fd_sc_hd__o2bb2ai_1 _19301_ (.A1_N(_08523_),
    .A2_N(_08544_),
    .B1(_08934_),
    .B2(_08936_),
    .Y(_08942_));
 sky130_fd_sc_hd__nand3_2 _19302_ (.A(_08942_),
    .B(net276),
    .C(_08941_),
    .Y(_08943_));
 sky130_fd_sc_hd__o211a_1 _19303_ (.A1(_08914_),
    .A2(net280),
    .B1(_04040_),
    .C1(_08925_),
    .X(_08944_));
 sky130_fd_sc_hd__o2bb2ai_2 _19304_ (.A1_N(_08935_),
    .A2_N(_08937_),
    .B1(_08938_),
    .B2(_08526_),
    .Y(_08945_));
 sky130_fd_sc_hd__o2111ai_4 _19305_ (.A1(_08521_),
    .A2(_02148_),
    .B1(_08937_),
    .C1(_08935_),
    .D1(_08939_),
    .Y(_08946_));
 sky130_fd_sc_hd__nand3_1 _19306_ (.A(_08945_),
    .B(_08946_),
    .C(net276),
    .Y(_08947_));
 sky130_fd_sc_hd__o31a_1 _19307_ (.A1(_04008_),
    .A2(net300),
    .A3(_08932_),
    .B1(_08947_),
    .X(_08948_));
 sky130_fd_sc_hd__a311o_1 _19308_ (.A1(_08945_),
    .A2(_08946_),
    .A3(net276),
    .B1(net273),
    .C1(_08944_),
    .X(_08949_));
 sky130_fd_sc_hd__o211ai_4 _19309_ (.A1(_02049_),
    .A2(net342),
    .B1(_08933_),
    .C1(_08943_),
    .Y(_08950_));
 sky130_fd_sc_hd__a311oi_4 _19310_ (.A1(_08945_),
    .A2(_08946_),
    .A3(net276),
    .B1(_08944_),
    .C1(_02148_),
    .Y(_08952_));
 sky130_fd_sc_hd__o211ai_4 _19311_ (.A1(net276),
    .A2(_08932_),
    .B1(_02137_),
    .C1(_08947_),
    .Y(_08953_));
 sky130_fd_sc_hd__a21oi_2 _19312_ (.A1(_08548_),
    .A2(net319),
    .B1(_08558_),
    .Y(_08954_));
 sky130_fd_sc_hd__o21ai_1 _19313_ (.A1(_08157_),
    .A2(_08556_),
    .B1(_08555_),
    .Y(_08955_));
 sky130_fd_sc_hd__o2bb2ai_4 _19314_ (.A1_N(_08555_),
    .A2_N(_08559_),
    .B1(_08542_),
    .B2(_08552_),
    .Y(_08956_));
 sky130_fd_sc_hd__o211ai_1 _19315_ (.A1(_08553_),
    .A2(_08954_),
    .B1(_08953_),
    .C1(_08950_),
    .Y(_08957_));
 sky130_fd_sc_hd__a21o_1 _19316_ (.A1(_08950_),
    .A2(_08953_),
    .B1(_08956_),
    .X(_08958_));
 sky130_fd_sc_hd__nand3_2 _19317_ (.A(_08958_),
    .B(net273),
    .C(_08957_),
    .Y(_08959_));
 sky130_fd_sc_hd__and3_1 _19318_ (.A(_05234_),
    .B(_08933_),
    .C(_08943_),
    .X(_08960_));
 sky130_fd_sc_hd__or2_2 _19319_ (.A(net273),
    .B(_08948_),
    .X(_08961_));
 sky130_fd_sc_hd__o2bb2ai_2 _19320_ (.A1_N(_08950_),
    .A2_N(_08953_),
    .B1(_08954_),
    .B2(_08553_),
    .Y(_08963_));
 sky130_fd_sc_hd__o2111ai_4 _19321_ (.A1(_08548_),
    .A2(net319),
    .B1(_08953_),
    .C1(_08950_),
    .D1(_08955_),
    .Y(_08964_));
 sky130_fd_sc_hd__nand3_2 _19322_ (.A(_08963_),
    .B(_08964_),
    .C(net273),
    .Y(_08965_));
 sky130_fd_sc_hd__and3_2 _19323_ (.A(_05486_),
    .B(_08949_),
    .C(_08959_),
    .X(_08966_));
 sky130_fd_sc_hd__a211o_2 _19324_ (.A1(_08961_),
    .A2(_08965_),
    .B1(_05481_),
    .C1(_05483_),
    .X(_08967_));
 sky130_fd_sc_hd__a311oi_4 _19325_ (.A1(_08963_),
    .A2(_08964_),
    .A3(net273),
    .B1(_08960_),
    .C1(net319),
    .Y(_08968_));
 sky130_fd_sc_hd__nand3_4 _19326_ (.A(_08965_),
    .B(net320),
    .C(_08961_),
    .Y(_08969_));
 sky130_fd_sc_hd__a22oi_1 _19327_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_08961_),
    .B2(_08965_),
    .Y(_08970_));
 sky130_fd_sc_hd__o211ai_4 _19328_ (.A1(_00174_),
    .A2(_00196_),
    .B1(_08949_),
    .C1(_08959_),
    .Y(_08971_));
 sky130_fd_sc_hd__o22a_1 _19329_ (.A1(_12888_),
    .A2(_08565_),
    .B1(_08569_),
    .B2(_08174_),
    .X(_08972_));
 sky130_fd_sc_hd__a21o_1 _19330_ (.A1(_08571_),
    .A2(_08573_),
    .B1(_08574_),
    .X(_08974_));
 sky130_fd_sc_hd__a21oi_2 _19331_ (.A1(_08573_),
    .A2(_08571_),
    .B1(_08574_),
    .Y(_08975_));
 sky130_fd_sc_hd__o2bb2ai_4 _19332_ (.A1_N(_08969_),
    .A2_N(_08971_),
    .B1(_08972_),
    .B2(_08572_),
    .Y(_08976_));
 sky130_fd_sc_hd__nand3_2 _19333_ (.A(_08974_),
    .B(_08971_),
    .C(_08969_),
    .Y(_08977_));
 sky130_fd_sc_hd__o311a_1 _19334_ (.A1(_08968_),
    .A2(_08970_),
    .A3(_08975_),
    .B1(net246),
    .C1(_08976_),
    .X(_08978_));
 sky130_fd_sc_hd__nand3_2 _19335_ (.A(_08976_),
    .B(_08977_),
    .C(net246),
    .Y(_08979_));
 sky130_fd_sc_hd__a31o_1 _19336_ (.A1(_08976_),
    .A2(_08977_),
    .A3(net246),
    .B1(_08966_),
    .X(_08980_));
 sky130_fd_sc_hd__and3_1 _19337_ (.A(_05754_),
    .B(_08967_),
    .C(_08979_),
    .X(_08981_));
 sky130_fd_sc_hd__a31oi_4 _19338_ (.A1(net330),
    .A2(_08567_),
    .A3(_08578_),
    .B1(_08591_),
    .Y(_08982_));
 sky130_fd_sc_hd__a22oi_4 _19339_ (.A1(_08190_),
    .A2(_08197_),
    .B1(_08584_),
    .B2(_11298_),
    .Y(_08983_));
 sky130_fd_sc_hd__a311oi_4 _19340_ (.A1(_08976_),
    .A2(_08977_),
    .A3(net246),
    .B1(_08966_),
    .C1(net326),
    .Y(_08985_));
 sky130_fd_sc_hd__a311o_2 _19341_ (.A1(_08976_),
    .A2(_08977_),
    .A3(net246),
    .B1(_08966_),
    .C1(net326),
    .X(_08986_));
 sky130_fd_sc_hd__a2bb2oi_4 _19342_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_08967_),
    .B2(_08979_),
    .Y(_08987_));
 sky130_fd_sc_hd__o22ai_4 _19343_ (.A1(net361),
    .A2(net345),
    .B1(_08966_),
    .B2(_08978_),
    .Y(_08988_));
 sky130_fd_sc_hd__o211ai_4 _19344_ (.A1(_08587_),
    .A2(_08982_),
    .B1(_08986_),
    .C1(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__o22ai_4 _19345_ (.A1(_08585_),
    .A2(_08983_),
    .B1(_08985_),
    .B2(_08987_),
    .Y(_08990_));
 sky130_fd_sc_hd__nand3_1 _19346_ (.A(_08989_),
    .B(_08990_),
    .C(net241),
    .Y(_08991_));
 sky130_fd_sc_hd__a21oi_2 _19347_ (.A1(_08967_),
    .A2(_08979_),
    .B1(net241),
    .Y(_08992_));
 sky130_fd_sc_hd__a211o_1 _19348_ (.A1(_08967_),
    .A2(_08979_),
    .B1(net266),
    .C1(_05751_),
    .X(_08993_));
 sky130_fd_sc_hd__o211ai_4 _19349_ (.A1(_08585_),
    .A2(_08983_),
    .B1(_08986_),
    .C1(_08988_),
    .Y(_08994_));
 sky130_fd_sc_hd__o22ai_4 _19350_ (.A1(_08587_),
    .A2(_08982_),
    .B1(_08985_),
    .B2(_08987_),
    .Y(_08996_));
 sky130_fd_sc_hd__o211ai_1 _19351_ (.A1(net266),
    .A2(_05751_),
    .B1(_08994_),
    .C1(_08996_),
    .Y(_08997_));
 sky130_fd_sc_hd__a31o_1 _19352_ (.A1(_08994_),
    .A2(_08996_),
    .A3(net241),
    .B1(_08992_),
    .X(_08998_));
 sky130_fd_sc_hd__a311oi_4 _19353_ (.A1(_08989_),
    .A2(_08990_),
    .A3(net241),
    .B1(_08981_),
    .C1(_11298_),
    .Y(_08999_));
 sky130_fd_sc_hd__o211ai_4 _19354_ (.A1(_08980_),
    .A2(net241),
    .B1(net330),
    .C1(_08991_),
    .Y(_09000_));
 sky130_fd_sc_hd__a311oi_4 _19355_ (.A1(_08994_),
    .A2(_08996_),
    .A3(net241),
    .B1(_08992_),
    .C1(_11309_),
    .Y(_09001_));
 sky130_fd_sc_hd__nand3_2 _19356_ (.A(_08997_),
    .B(_11298_),
    .C(_08993_),
    .Y(_09002_));
 sky130_fd_sc_hd__a21oi_1 _19357_ (.A1(net348),
    .A2(_08598_),
    .B1(_08607_),
    .Y(_09003_));
 sky130_fd_sc_hd__o2111ai_1 _19358_ (.A1(_10015_),
    .A2(_08597_),
    .B1(_08610_),
    .C1(_09000_),
    .D1(_09002_),
    .Y(_09004_));
 sky130_fd_sc_hd__o22ai_1 _19359_ (.A1(_08600_),
    .A2(_08609_),
    .B1(_08999_),
    .B2(_09001_),
    .Y(_09005_));
 sky130_fd_sc_hd__o211ai_2 _19360_ (.A1(net259),
    .A2(net257),
    .B1(_09004_),
    .C1(_09005_),
    .Y(_09007_));
 sky130_fd_sc_hd__a311o_4 _19361_ (.A1(_08989_),
    .A2(_08990_),
    .A3(net241),
    .B1(net240),
    .C1(_08981_),
    .X(_09008_));
 sky130_fd_sc_hd__o2bb2ai_1 _19362_ (.A1_N(_09000_),
    .A2_N(_09002_),
    .B1(_09003_),
    .B2(_08603_),
    .Y(_09009_));
 sky130_fd_sc_hd__o21ai_1 _19363_ (.A1(_08600_),
    .A2(_08609_),
    .B1(_09000_),
    .Y(_09010_));
 sky130_fd_sc_hd__o221ai_4 _19364_ (.A1(net259),
    .A2(net257),
    .B1(_09001_),
    .B2(_09010_),
    .C1(_09009_),
    .Y(_09011_));
 sky130_fd_sc_hd__nand2_1 _19365_ (.A(_09008_),
    .B(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__and3_1 _19366_ (.A(_06294_),
    .B(_09008_),
    .C(_09011_),
    .X(_09013_));
 sky130_fd_sc_hd__or3_2 _19367_ (.A(_06291_),
    .B(_06292_),
    .C(_09012_),
    .X(_09014_));
 sky130_fd_sc_hd__a2bb2oi_2 _19368_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_09008_),
    .B2(_09011_),
    .Y(_09015_));
 sky130_fd_sc_hd__o211ai_4 _19369_ (.A1(_08998_),
    .A2(net240),
    .B1(_10025_),
    .C1(_09007_),
    .Y(_09016_));
 sky130_fd_sc_hd__o211a_2 _19370_ (.A1(net365),
    .A2(net364),
    .B1(_09008_),
    .C1(_09011_),
    .X(_09018_));
 sky130_fd_sc_hd__o211ai_4 _19371_ (.A1(net365),
    .A2(net364),
    .B1(_09008_),
    .C1(_09011_),
    .Y(_09019_));
 sky130_fd_sc_hd__o21a_1 _19372_ (.A1(_08224_),
    .A2(_08231_),
    .B1(_08619_),
    .X(_09020_));
 sky130_fd_sc_hd__o21ai_2 _19373_ (.A1(_08224_),
    .A2(_08231_),
    .B1(_08619_),
    .Y(_09021_));
 sky130_fd_sc_hd__a21oi_2 _19374_ (.A1(_08619_),
    .A2(_08624_),
    .B1(_08620_),
    .Y(_09022_));
 sky130_fd_sc_hd__o2bb2ai_1 _19375_ (.A1_N(_09016_),
    .A2_N(_09019_),
    .B1(_09020_),
    .B2(_08620_),
    .Y(_09023_));
 sky130_fd_sc_hd__nand4_2 _19376_ (.A(_08621_),
    .B(_09016_),
    .C(_09019_),
    .D(_09021_),
    .Y(_09024_));
 sky130_fd_sc_hd__nand3_2 _19377_ (.A(_09023_),
    .B(_09024_),
    .C(net212),
    .Y(_09025_));
 sky130_fd_sc_hd__a22o_1 _19378_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_09008_),
    .B2(_09011_),
    .X(_09026_));
 sky130_fd_sc_hd__o21ai_1 _19379_ (.A1(_09015_),
    .A2(_09018_),
    .B1(_09022_),
    .Y(_09027_));
 sky130_fd_sc_hd__o22a_1 _19380_ (.A1(_10025_),
    .A2(_09012_),
    .B1(_09020_),
    .B2(_08620_),
    .X(_09029_));
 sky130_fd_sc_hd__o211ai_1 _19381_ (.A1(_08620_),
    .A2(_09020_),
    .B1(_09019_),
    .C1(_09016_),
    .Y(_09030_));
 sky130_fd_sc_hd__nand3_1 _19382_ (.A(_09027_),
    .B(_09030_),
    .C(net212),
    .Y(_09031_));
 sky130_fd_sc_hd__a31o_1 _19383_ (.A1(_09023_),
    .A2(_09024_),
    .A3(net212),
    .B1(_09013_),
    .X(_09032_));
 sky130_fd_sc_hd__nand3_2 _19384_ (.A(_09031_),
    .B(_08907_),
    .C(_09026_),
    .Y(_09033_));
 sky130_fd_sc_hd__and3_1 _19385_ (.A(_08918_),
    .B(_09014_),
    .C(_09025_),
    .X(_09034_));
 sky130_fd_sc_hd__o211ai_1 _19386_ (.A1(_08819_),
    .A2(_08841_),
    .B1(_09014_),
    .C1(_09025_),
    .Y(_09035_));
 sky130_fd_sc_hd__nand3_1 _19387_ (.A(_08722_),
    .B(_09033_),
    .C(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__a21o_1 _19388_ (.A1(_09033_),
    .A2(_09035_),
    .B1(_08722_),
    .X(_09037_));
 sky130_fd_sc_hd__nand3_2 _19389_ (.A(_09037_),
    .B(net211),
    .C(_09036_),
    .Y(_09038_));
 sky130_fd_sc_hd__a311o_1 _19390_ (.A1(_09023_),
    .A2(_09024_),
    .A3(net212),
    .B1(net211),
    .C1(_09013_),
    .X(_09040_));
 sky130_fd_sc_hd__o31a_1 _19391_ (.A1(_06608_),
    .A2(net237),
    .A3(_09032_),
    .B1(_09038_),
    .X(_09041_));
 sky130_fd_sc_hd__inv_2 _19392_ (.A(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__a22oi_2 _19393_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_09038_),
    .B2(_09040_),
    .Y(_09043_));
 sky130_fd_sc_hd__a22o_1 _19394_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_09038_),
    .B2(_09040_),
    .X(_09044_));
 sky130_fd_sc_hd__o221a_1 _19395_ (.A1(net368),
    .A2(_07866_),
    .B1(net211),
    .B2(_09032_),
    .C1(_09038_),
    .X(_09045_));
 sky130_fd_sc_hd__o221ai_4 _19396_ (.A1(net368),
    .A2(_07866_),
    .B1(net211),
    .B2(_09032_),
    .C1(_09038_),
    .Y(_09046_));
 sky130_fd_sc_hd__a32oi_4 _19397_ (.A1(_08644_),
    .A2(_06978_),
    .A3(_06956_),
    .B1(_08651_),
    .B2(_08648_),
    .Y(_09047_));
 sky130_fd_sc_hd__a21boi_2 _19398_ (.A1(_08649_),
    .A2(_08650_),
    .B1_N(_08651_),
    .Y(_09048_));
 sky130_fd_sc_hd__o21ai_1 _19399_ (.A1(_09043_),
    .A2(_09045_),
    .B1(_09047_),
    .Y(_09049_));
 sky130_fd_sc_hd__nand3_1 _19400_ (.A(_09044_),
    .B(_09046_),
    .C(_09048_),
    .Y(_09051_));
 sky130_fd_sc_hd__o21ai_1 _19401_ (.A1(_09043_),
    .A2(_09045_),
    .B1(_09048_),
    .Y(_09052_));
 sky130_fd_sc_hd__nand2_1 _19402_ (.A(_09047_),
    .B(_09046_),
    .Y(_09053_));
 sky130_fd_sc_hd__o221ai_1 _19403_ (.A1(net230),
    .A2(_06901_),
    .B1(_09043_),
    .B2(_09053_),
    .C1(_09052_),
    .Y(_09054_));
 sky130_fd_sc_hd__nand3_4 _19404_ (.A(_09049_),
    .B(_09051_),
    .C(net208),
    .Y(_09055_));
 sky130_fd_sc_hd__o21ai_2 _19405_ (.A1(_06897_),
    .A2(_06898_),
    .B1(_09041_),
    .Y(_09056_));
 sky130_fd_sc_hd__o21ai_2 _19406_ (.A1(net208),
    .A2(_09042_),
    .B1(_09055_),
    .Y(_09057_));
 sky130_fd_sc_hd__and3_1 _19407_ (.A(_09055_),
    .B(_09056_),
    .C(_07232_),
    .X(_09058_));
 sky130_fd_sc_hd__or3_1 _19408_ (.A(_07227_),
    .B(net203),
    .C(_09057_),
    .X(_09059_));
 sky130_fd_sc_hd__a31oi_1 _19409_ (.A1(_08658_),
    .A2(_06332_),
    .A3(_08647_),
    .B1(_08664_),
    .Y(_09060_));
 sky130_fd_sc_hd__nor2_1 _19410_ (.A(_08665_),
    .B(_08662_),
    .Y(_09062_));
 sky130_fd_sc_hd__o21ai_1 _19411_ (.A1(_08665_),
    .A2(_08662_),
    .B1(_08661_),
    .Y(_09063_));
 sky130_fd_sc_hd__a22oi_4 _19412_ (.A1(net376),
    .A2(_07022_),
    .B1(_09055_),
    .B2(_09056_),
    .Y(_09064_));
 sky130_fd_sc_hd__o221ai_1 _19413_ (.A1(_06989_),
    .A2(net375),
    .B1(net208),
    .B2(_09041_),
    .C1(_09054_),
    .Y(_09065_));
 sky130_fd_sc_hd__o211a_1 _19414_ (.A1(_09042_),
    .A2(net208),
    .B1(_07044_),
    .C1(_09055_),
    .X(_09066_));
 sky130_fd_sc_hd__o211ai_2 _19415_ (.A1(_09042_),
    .A2(net208),
    .B1(_07044_),
    .C1(_09055_),
    .Y(_09067_));
 sky130_fd_sc_hd__o21ai_2 _19416_ (.A1(_08662_),
    .A2(_09060_),
    .B1(_09067_),
    .Y(_09068_));
 sky130_fd_sc_hd__o22ai_2 _19417_ (.A1(_08660_),
    .A2(_09062_),
    .B1(_09064_),
    .B2(_09066_),
    .Y(_09069_));
 sky130_fd_sc_hd__o211a_1 _19418_ (.A1(_09068_),
    .A2(_09064_),
    .B1(net185),
    .C1(_09069_),
    .X(_09070_));
 sky130_fd_sc_hd__o211ai_4 _19419_ (.A1(_09068_),
    .A2(_09064_),
    .B1(net185),
    .C1(_09069_),
    .Y(_09071_));
 sky130_fd_sc_hd__o31a_1 _19420_ (.A1(_07227_),
    .A2(net203),
    .A3(_09057_),
    .B1(_09071_),
    .X(_09073_));
 sky130_fd_sc_hd__or3_1 _19421_ (.A(_07544_),
    .B(net184),
    .C(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__a2bb2oi_2 _19422_ (.A1_N(net394),
    .A2_N(_06267_),
    .B1(_09059_),
    .B2(_09071_),
    .Y(_09075_));
 sky130_fd_sc_hd__a22o_1 _19423_ (.A1(_06256_),
    .A2(_06278_),
    .B1(_09059_),
    .B2(_09071_),
    .X(_09076_));
 sky130_fd_sc_hd__o21ai_1 _19424_ (.A1(net381),
    .A2(_06310_),
    .B1(_09071_),
    .Y(_09077_));
 sky130_fd_sc_hd__o221a_1 _19425_ (.A1(net381),
    .A2(_06310_),
    .B1(net185),
    .B2(_09057_),
    .C1(_09071_),
    .X(_09078_));
 sky130_fd_sc_hd__a31oi_1 _19426_ (.A1(_08659_),
    .A2(_08669_),
    .A3(_08672_),
    .B1(_08671_),
    .Y(_09079_));
 sky130_fd_sc_hd__a31o_1 _19427_ (.A1(_08659_),
    .A2(_08669_),
    .A3(_08672_),
    .B1(_08671_),
    .X(_09080_));
 sky130_fd_sc_hd__o21ai_1 _19428_ (.A1(_09075_),
    .A2(_09078_),
    .B1(_09079_),
    .Y(_09081_));
 sky130_fd_sc_hd__o211ai_1 _19429_ (.A1(_09058_),
    .A2(_09077_),
    .B1(_09080_),
    .C1(_09076_),
    .Y(_09082_));
 sky130_fd_sc_hd__o21ai_1 _19430_ (.A1(_09075_),
    .A2(_09078_),
    .B1(_09080_),
    .Y(_09084_));
 sky130_fd_sc_hd__o31a_1 _19431_ (.A1(_06343_),
    .A2(_09058_),
    .A3(_09070_),
    .B1(_09079_),
    .X(_09085_));
 sky130_fd_sc_hd__a31o_2 _19432_ (.A1(_06332_),
    .A2(_09059_),
    .A3(_09071_),
    .B1(_09080_),
    .X(_09086_));
 sky130_fd_sc_hd__o221ai_4 _19433_ (.A1(_07544_),
    .A2(net184),
    .B1(_09075_),
    .B2(_09086_),
    .C1(_09084_),
    .Y(_09087_));
 sky130_fd_sc_hd__o211a_1 _19434_ (.A1(_07544_),
    .A2(net184),
    .B1(_09081_),
    .C1(_09082_),
    .X(_09088_));
 sky130_fd_sc_hd__o311a_1 _19435_ (.A1(_07227_),
    .A2(net203),
    .A3(_09057_),
    .B1(_09071_),
    .C1(_07550_),
    .X(_09089_));
 sky130_fd_sc_hd__a22oi_1 _19436_ (.A1(_05545_),
    .A2(_08680_),
    .B1(_08676_),
    .B2(_08675_),
    .Y(_09090_));
 sky130_fd_sc_hd__a22o_1 _19437_ (.A1(_05545_),
    .A2(_08680_),
    .B1(_08676_),
    .B2(_08675_),
    .X(_09091_));
 sky130_fd_sc_hd__and3_1 _19438_ (.A(_09091_),
    .B(_05851_),
    .C(_08682_),
    .X(_09092_));
 sky130_fd_sc_hd__o211ai_2 _19439_ (.A1(_05545_),
    .A2(_08680_),
    .B1(_05851_),
    .C1(_09091_),
    .Y(_09093_));
 sky130_fd_sc_hd__o21ai_2 _19440_ (.A1(_08681_),
    .A2(_09090_),
    .B1(_05862_),
    .Y(_09095_));
 sky130_fd_sc_hd__o211ai_4 _19441_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_09093_),
    .C1(_09095_),
    .Y(_09096_));
 sky130_fd_sc_hd__o211a_1 _19442_ (.A1(net163),
    .A2(_09073_),
    .B1(_09087_),
    .C1(_09096_),
    .X(_09097_));
 sky130_fd_sc_hd__o211ai_2 _19443_ (.A1(net163),
    .A2(_09073_),
    .B1(_09087_),
    .C1(_09096_),
    .Y(_09098_));
 sky130_fd_sc_hd__a21oi_2 _19444_ (.A1(_09074_),
    .A2(_09087_),
    .B1(_09096_),
    .Y(_09099_));
 sky130_fd_sc_hd__o31a_1 _19445_ (.A1(_09096_),
    .A2(_09089_),
    .A3(_09088_),
    .B1(_09098_),
    .X(_09100_));
 sky130_fd_sc_hd__o32ai_1 _19446_ (.A1(_05250_),
    .A2(_08686_),
    .A3(_08688_),
    .B1(_08290_),
    .B2(_08696_),
    .Y(_09101_));
 sky130_fd_sc_hd__o221ai_4 _19447_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_08290_),
    .B2(_08696_),
    .C1(_08695_),
    .Y(_09102_));
 sky130_fd_sc_hd__o22ai_4 _19448_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_08694_),
    .B2(_08698_),
    .Y(_09103_));
 sky130_fd_sc_hd__a22oi_1 _19449_ (.A1(_08297_),
    .A2(_08299_),
    .B1(_09101_),
    .B2(_05556_),
    .Y(_09104_));
 sky130_fd_sc_hd__o211ai_2 _19450_ (.A1(net180),
    .A2(_08298_),
    .B1(_09102_),
    .C1(_09103_),
    .Y(_09106_));
 sky130_fd_sc_hd__nor3_1 _19451_ (.A(_09097_),
    .B(_09099_),
    .C(_09106_),
    .Y(_09107_));
 sky130_fd_sc_hd__nand3_1 _19452_ (.A(_09100_),
    .B(_09102_),
    .C(_09104_),
    .Y(_09108_));
 sky130_fd_sc_hd__a21oi_1 _19453_ (.A1(_09104_),
    .A2(_09102_),
    .B1(_09100_),
    .Y(_09109_));
 sky130_fd_sc_hd__o21ai_2 _19454_ (.A1(_09097_),
    .A2(_09099_),
    .B1(_09106_),
    .Y(_09110_));
 sky130_fd_sc_hd__o31a_1 _19455_ (.A1(_09097_),
    .A2(_09099_),
    .A3(_09106_),
    .B1(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__o311a_1 _19456_ (.A1(_09097_),
    .A2(_09099_),
    .A3(_09106_),
    .B1(_05239_),
    .C1(_09110_),
    .X(_09112_));
 sky130_fd_sc_hd__a21oi_2 _19457_ (.A1(_09108_),
    .A2(_09110_),
    .B1(_05239_),
    .Y(_09113_));
 sky130_fd_sc_hd__o21ai_1 _19458_ (.A1(_09112_),
    .A2(_09113_),
    .B1(_08702_),
    .Y(_09114_));
 sky130_fd_sc_hd__o31a_1 _19459_ (.A1(_08702_),
    .A2(_09112_),
    .A3(_09113_),
    .B1(_08714_),
    .X(_09115_));
 sky130_fd_sc_hd__a22oi_2 _19460_ (.A1(_08715_),
    .A2(_09111_),
    .B1(_09115_),
    .B2(_09114_),
    .Y(_09117_));
 sky130_fd_sc_hd__or3_4 _19461_ (.A(net48),
    .B(net49),
    .C(_08292_),
    .X(_09118_));
 sky130_fd_sc_hd__o21ai_4 _19462_ (.A1(net49),
    .A2(_08704_),
    .B1(net409),
    .Y(_09119_));
 sky130_fd_sc_hd__nor2_8 _19463_ (.A(net50),
    .B(_09119_),
    .Y(_09120_));
 sky130_fd_sc_hd__and2_4 _19464_ (.A(_09119_),
    .B(net50),
    .X(_09121_));
 sky130_fd_sc_hd__o311a_4 _19465_ (.A1(net48),
    .A2(net49),
    .A3(_08292_),
    .B1(net50),
    .C1(net409),
    .X(_09122_));
 sky130_fd_sc_hd__a21oi_4 _19466_ (.A1(_09118_),
    .A2(net409),
    .B1(net50),
    .Y(_09123_));
 sky130_fd_sc_hd__or2_4 _19467_ (.A(_09122_),
    .B(_09123_),
    .X(_09124_));
 sky130_fd_sc_hd__nor2_8 _19468_ (.A(_09122_),
    .B(_09123_),
    .Y(_09125_));
 sky130_fd_sc_hd__o21ai_1 _19469_ (.A1(_03289_),
    .A2(_09124_),
    .B1(_09117_),
    .Y(_09126_));
 sky130_fd_sc_hd__nor2_1 _19470_ (.A(_03289_),
    .B(_09117_),
    .Y(_09128_));
 sky130_fd_sc_hd__o31ai_1 _19471_ (.A1(_03289_),
    .A2(_09117_),
    .A3(_09124_),
    .B1(_09126_),
    .Y(_09129_));
 sky130_fd_sc_hd__xnor2_1 _19472_ (.A(_08720_),
    .B(_09129_),
    .Y(net82));
 sky130_fd_sc_hd__and3_1 _19473_ (.A(_09129_),
    .B(_08717_),
    .C(_08305_),
    .X(_09130_));
 sky130_fd_sc_hd__a21oi_1 _19474_ (.A1(_09047_),
    .A2(_09046_),
    .B1(_09043_),
    .Y(_09131_));
 sky130_fd_sc_hd__o21ai_2 _19475_ (.A1(_09048_),
    .A2(_09045_),
    .B1(_09044_),
    .Y(_09132_));
 sky130_fd_sc_hd__or4_4 _19476_ (.A(net16),
    .B(net17),
    .C(net18),
    .D(_07926_),
    .X(_09133_));
 sky130_fd_sc_hd__and3b_4 _19477_ (.A_N(net19),
    .B(_09133_),
    .C(net410),
    .X(_09134_));
 sky130_fd_sc_hd__a21boi_4 _19478_ (.A1(_09133_),
    .A2(net410),
    .B1_N(net19),
    .Y(_09135_));
 sky130_fd_sc_hd__o311a_4 _19479_ (.A1(net17),
    .A2(net18),
    .A3(_08306_),
    .B1(net19),
    .C1(net410),
    .X(_09136_));
 sky130_fd_sc_hd__a21oi_4 _19480_ (.A1(_09133_),
    .A2(net410),
    .B1(net19),
    .Y(_09138_));
 sky130_fd_sc_hd__nor2_8 _19481_ (.A(net194),
    .B(net191),
    .Y(_09139_));
 sky130_fd_sc_hd__nor2_8 _19482_ (.A(_09136_),
    .B(_09138_),
    .Y(_09140_));
 sky130_fd_sc_hd__o21a_1 _19483_ (.A1(_09134_),
    .A2(_09135_),
    .B1(net33),
    .X(_09141_));
 sky130_fd_sc_hd__or3_2 _19484_ (.A(_03178_),
    .B(_09136_),
    .C(_09138_),
    .X(_09142_));
 sky130_fd_sc_hd__a22oi_4 _19485_ (.A1(_08316_),
    .A2(net175),
    .B1(_08739_),
    .B2(_08744_),
    .Y(_09143_));
 sky130_fd_sc_hd__or3_1 _19486_ (.A(_08724_),
    .B(_08726_),
    .C(_09141_),
    .X(_09144_));
 sky130_fd_sc_hd__o21ai_4 _19487_ (.A1(_08733_),
    .A2(net174),
    .B1(_09144_),
    .Y(_09145_));
 sky130_fd_sc_hd__a21oi_2 _19488_ (.A1(_08742_),
    .A2(_08747_),
    .B1(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__o311a_1 _19489_ (.A1(_08311_),
    .A2(_08733_),
    .A3(_08312_),
    .B1(_09145_),
    .C1(_08747_),
    .X(_09147_));
 sky130_fd_sc_hd__a31o_1 _19490_ (.A1(_08742_),
    .A2(_08747_),
    .A3(_09145_),
    .B1(_05185_),
    .X(_09149_));
 sky130_fd_sc_hd__o32a_1 _19491_ (.A1(_03178_),
    .A2(_09136_),
    .A3(_09138_),
    .B1(_05130_),
    .B2(_05152_),
    .X(_09150_));
 sky130_fd_sc_hd__o211a_1 _19492_ (.A1(_09146_),
    .A2(_09147_),
    .B1(_05141_),
    .C1(_05163_),
    .X(_09151_));
 sky130_fd_sc_hd__o22ai_4 _19493_ (.A1(net405),
    .A2(_09142_),
    .B1(_09146_),
    .B2(_09149_),
    .Y(_09152_));
 sky130_fd_sc_hd__inv_2 _19494_ (.A(_09152_),
    .Y(_09153_));
 sky130_fd_sc_hd__and3_1 _19495_ (.A(_05359_),
    .B(_05381_),
    .C(_09152_),
    .X(_09154_));
 sky130_fd_sc_hd__or4_1 _19496_ (.A(_05348_),
    .B(net401),
    .C(_09150_),
    .D(_09151_),
    .X(_09155_));
 sky130_fd_sc_hd__o21a_1 _19497_ (.A1(_08307_),
    .A2(_08309_),
    .B1(_09152_),
    .X(_09156_));
 sky130_fd_sc_hd__or4_1 _19498_ (.A(_08311_),
    .B(_08312_),
    .C(_09150_),
    .D(_09151_),
    .X(_09157_));
 sky130_fd_sc_hd__o221a_1 _19499_ (.A1(net405),
    .A2(_09142_),
    .B1(_09146_),
    .B2(_09149_),
    .C1(net199),
    .X(_09158_));
 sky130_fd_sc_hd__nor2_1 _19500_ (.A(_09156_),
    .B(_09158_),
    .Y(_09160_));
 sky130_fd_sc_hd__nand4_2 _19501_ (.A(_08333_),
    .B(_07954_),
    .C(_07584_),
    .D(_08330_),
    .Y(_09161_));
 sky130_fd_sc_hd__and4b_2 _19502_ (.A_N(_09161_),
    .B(_08753_),
    .C(_08751_),
    .D(_07594_),
    .X(_09162_));
 sky130_fd_sc_hd__nand4b_2 _19503_ (.A_N(_09161_),
    .B(_08753_),
    .C(_08751_),
    .D(_07594_),
    .Y(_09163_));
 sky130_fd_sc_hd__o21ai_2 _19504_ (.A1(_08750_),
    .A2(_09161_),
    .B1(_08753_),
    .Y(_09164_));
 sky130_fd_sc_hd__a21oi_4 _19505_ (.A1(_08758_),
    .A2(_08755_),
    .B1(_09164_),
    .Y(_09165_));
 sky130_fd_sc_hd__o21bai_2 _19506_ (.A1(_08756_),
    .A2(_08757_),
    .B1_N(_09164_),
    .Y(_09166_));
 sky130_fd_sc_hd__nor2_1 _19507_ (.A(_09162_),
    .B(_09165_),
    .Y(_09167_));
 sky130_fd_sc_hd__nand3_2 _19508_ (.A(_09166_),
    .B(_09160_),
    .C(_09163_),
    .Y(_09168_));
 sky130_fd_sc_hd__o22ai_4 _19509_ (.A1(_09156_),
    .A2(_09158_),
    .B1(_09162_),
    .B2(_09165_),
    .Y(_09169_));
 sky130_fd_sc_hd__o211a_1 _19510_ (.A1(_05348_),
    .A2(net401),
    .B1(_09168_),
    .C1(_09169_),
    .X(_09171_));
 sky130_fd_sc_hd__o211ai_4 _19511_ (.A1(_05348_),
    .A2(net401),
    .B1(_09168_),
    .C1(_09169_),
    .Y(_09172_));
 sky130_fd_sc_hd__o31a_1 _19512_ (.A1(_05403_),
    .A2(_09150_),
    .A3(_09151_),
    .B1(_09172_),
    .X(_09173_));
 sky130_fd_sc_hd__a31o_1 _19513_ (.A1(_05403_),
    .A2(_09168_),
    .A3(_09169_),
    .B1(_09154_),
    .X(_09174_));
 sky130_fd_sc_hd__and3_1 _19514_ (.A(_05687_),
    .B(_05709_),
    .C(_09174_),
    .X(_09175_));
 sky130_fd_sc_hd__or3_1 _19515_ (.A(_05676_),
    .B(_05698_),
    .C(_09173_),
    .X(_09176_));
 sky130_fd_sc_hd__a2bb2oi_2 _19516_ (.A1_N(_07928_),
    .A2_N(_07930_),
    .B1(_09155_),
    .B2(_09172_),
    .Y(_09177_));
 sky130_fd_sc_hd__o22ai_4 _19517_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_09154_),
    .B2(_09171_),
    .Y(_09178_));
 sky130_fd_sc_hd__a31oi_1 _19518_ (.A1(_05403_),
    .A2(_09168_),
    .A3(_09169_),
    .B1(_07936_),
    .Y(_09179_));
 sky130_fd_sc_hd__o311a_1 _19519_ (.A1(_05403_),
    .A2(_09150_),
    .A3(_09151_),
    .B1(_07935_),
    .C1(_09172_),
    .X(_09180_));
 sky130_fd_sc_hd__o211ai_4 _19520_ (.A1(_05403_),
    .A2(_09153_),
    .B1(_07935_),
    .C1(_09172_),
    .Y(_09182_));
 sky130_fd_sc_hd__a21oi_2 _19521_ (.A1(_09155_),
    .A2(_09179_),
    .B1(_09177_),
    .Y(_09183_));
 sky130_fd_sc_hd__nand2_1 _19522_ (.A(_09178_),
    .B(_09182_),
    .Y(_09184_));
 sky130_fd_sc_hd__a21oi_1 _19523_ (.A1(_08773_),
    .A2(_08770_),
    .B1(_08767_),
    .Y(_09185_));
 sky130_fd_sc_hd__o32ai_4 _19524_ (.A1(_07564_),
    .A2(_08762_),
    .A3(_08763_),
    .B1(_08771_),
    .B2(_08772_),
    .Y(_09186_));
 sky130_fd_sc_hd__nand2_2 _19525_ (.A(_09186_),
    .B(_09183_),
    .Y(_09187_));
 sky130_fd_sc_hd__o221ai_4 _19526_ (.A1(_08771_),
    .A2(_08772_),
    .B1(_09177_),
    .B2(_09180_),
    .C1(_08768_),
    .Y(_09188_));
 sky130_fd_sc_hd__nand3_1 _19527_ (.A(_09187_),
    .B(_09188_),
    .C(net358),
    .Y(_09189_));
 sky130_fd_sc_hd__a22o_1 _19528_ (.A1(_05687_),
    .A2(_05709_),
    .B1(_09187_),
    .B2(_09188_),
    .X(_09190_));
 sky130_fd_sc_hd__o31a_2 _19529_ (.A1(_05676_),
    .A2(_05698_),
    .A3(_09173_),
    .B1(_09189_),
    .X(_09191_));
 sky130_fd_sc_hd__a2bb2oi_2 _19530_ (.A1_N(_07555_),
    .A2_N(net218),
    .B1(_09176_),
    .B2(_09189_),
    .Y(_09193_));
 sky130_fd_sc_hd__a22o_1 _19531_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_09176_),
    .B2(_09189_),
    .X(_09194_));
 sky130_fd_sc_hd__a311oi_4 _19532_ (.A1(_09187_),
    .A2(_09188_),
    .A3(net358),
    .B1(net202),
    .C1(_09175_),
    .Y(_09195_));
 sky130_fd_sc_hd__a311o_2 _19533_ (.A1(_09187_),
    .A2(_09188_),
    .A3(net358),
    .B1(net202),
    .C1(_09175_),
    .X(_09196_));
 sky130_fd_sc_hd__nor2_1 _19534_ (.A(_09193_),
    .B(_09195_),
    .Y(_09197_));
 sky130_fd_sc_hd__nand2_1 _19535_ (.A(_09194_),
    .B(_09196_),
    .Y(_09198_));
 sky130_fd_sc_hd__a21oi_1 _19536_ (.A1(_08791_),
    .A2(_08788_),
    .B1(_08784_),
    .Y(_09199_));
 sky130_fd_sc_hd__o32ai_1 _19537_ (.A1(_07244_),
    .A2(_07245_),
    .A3(_08780_),
    .B1(_08789_),
    .B2(_08790_),
    .Y(_09200_));
 sky130_fd_sc_hd__o221a_1 _19538_ (.A1(_09193_),
    .A2(_09195_),
    .B1(_08789_),
    .B2(_08790_),
    .C1(_08785_),
    .X(_09201_));
 sky130_fd_sc_hd__o221ai_4 _19539_ (.A1(_08789_),
    .A2(_08790_),
    .B1(_09193_),
    .B2(_09195_),
    .C1(_08785_),
    .Y(_09202_));
 sky130_fd_sc_hd__nand2_2 _19540_ (.A(_09200_),
    .B(_09197_),
    .Y(_09204_));
 sky130_fd_sc_hd__o311a_2 _19541_ (.A1(_05676_),
    .A2(_09174_),
    .A3(_05698_),
    .B1(_06848_),
    .C1(_09190_),
    .X(_09205_));
 sky130_fd_sc_hd__or3_1 _19542_ (.A(_06793_),
    .B(_06815_),
    .C(_09191_),
    .X(_09206_));
 sky130_fd_sc_hd__o22ai_2 _19543_ (.A1(net379),
    .A2(net378),
    .B1(_09198_),
    .B2(_09199_),
    .Y(_09207_));
 sky130_fd_sc_hd__nand3_1 _19544_ (.A(_09204_),
    .B(net357),
    .C(_09202_),
    .Y(_09208_));
 sky130_fd_sc_hd__o22ai_2 _19545_ (.A1(net357),
    .A2(_09191_),
    .B1(_09201_),
    .B2(_09207_),
    .Y(_09209_));
 sky130_fd_sc_hd__o22a_4 _19546_ (.A1(net357),
    .A2(_09191_),
    .B1(_09201_),
    .B2(_09207_),
    .X(_09210_));
 sky130_fd_sc_hd__or3_1 _19547_ (.A(_07691_),
    .B(net371),
    .C(_09210_),
    .X(_09211_));
 sky130_fd_sc_hd__a2bb2oi_1 _19548_ (.A1_N(_07242_),
    .A2_N(_07243_),
    .B1(_09206_),
    .B2(_09208_),
    .Y(_09212_));
 sky130_fd_sc_hd__o21ai_4 _19549_ (.A1(_07242_),
    .A2(_07243_),
    .B1(_09209_),
    .Y(_09213_));
 sky130_fd_sc_hd__a31o_1 _19550_ (.A1(_09204_),
    .A2(net357),
    .A3(_09202_),
    .B1(net222),
    .X(_09215_));
 sky130_fd_sc_hd__a311oi_4 _19551_ (.A1(_09204_),
    .A2(net357),
    .A3(_09202_),
    .B1(_09205_),
    .C1(net222),
    .Y(_09216_));
 sky130_fd_sc_hd__a311o_1 _19552_ (.A1(_09204_),
    .A2(net357),
    .A3(_09202_),
    .B1(_09205_),
    .C1(net222),
    .X(_09217_));
 sky130_fd_sc_hd__a2bb2oi_1 _19553_ (.A1_N(net227),
    .A2_N(_08798_),
    .B1(_08811_),
    .B2(_08813_),
    .Y(_09218_));
 sky130_fd_sc_hd__o22ai_2 _19554_ (.A1(net227),
    .A2(_08798_),
    .B1(_08810_),
    .B2(_08812_),
    .Y(_09219_));
 sky130_fd_sc_hd__o211ai_1 _19555_ (.A1(net225),
    .A2(_08799_),
    .B1(_08811_),
    .C1(_08813_),
    .Y(_09220_));
 sky130_fd_sc_hd__o21ai_1 _19556_ (.A1(net227),
    .A2(_08798_),
    .B1(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__o2111ai_4 _19557_ (.A1(net225),
    .A2(_08799_),
    .B1(_09213_),
    .C1(_09217_),
    .D1(_09219_),
    .Y(_09222_));
 sky130_fd_sc_hd__o211ai_2 _19558_ (.A1(_09212_),
    .A2(_09216_),
    .B1(_08801_),
    .C1(_08816_),
    .Y(_09223_));
 sky130_fd_sc_hd__nand3_4 _19559_ (.A(_09223_),
    .B(net355),
    .C(_09222_),
    .Y(_09224_));
 sky130_fd_sc_hd__o31a_1 _19560_ (.A1(net374),
    .A2(_07702_),
    .A3(_09210_),
    .B1(_09224_),
    .X(_09226_));
 sky130_fd_sc_hd__o21ai_2 _19561_ (.A1(net354),
    .A2(_09210_),
    .B1(_09224_),
    .Y(_09227_));
 sky130_fd_sc_hd__a2bb2oi_2 _19562_ (.A1_N(_06914_),
    .A2_N(_06916_),
    .B1(_09211_),
    .B2(_09224_),
    .Y(_09228_));
 sky130_fd_sc_hd__a22o_2 _19563_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_09211_),
    .B2(_09224_),
    .X(_09229_));
 sky130_fd_sc_hd__o221a_1 _19564_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_09210_),
    .B2(net354),
    .C1(_09224_),
    .X(_09230_));
 sky130_fd_sc_hd__o221ai_4 _19565_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_09210_),
    .B2(net354),
    .C1(_09224_),
    .Y(_09231_));
 sky130_fd_sc_hd__nor2_1 _19566_ (.A(_09228_),
    .B(_09230_),
    .Y(_09232_));
 sky130_fd_sc_hd__o211a_1 _19567_ (.A1(_08022_),
    .A2(_08028_),
    .B1(_07655_),
    .C1(_08027_),
    .X(_09233_));
 sky130_fd_sc_hd__nand4_1 _19568_ (.A(_08412_),
    .B(_09233_),
    .C(_08417_),
    .D(_07664_),
    .Y(_09234_));
 sky130_fd_sc_hd__nor3_2 _19569_ (.A(_09234_),
    .B(_08831_),
    .C(_08828_),
    .Y(_09235_));
 sky130_fd_sc_hd__nand3b_2 _19570_ (.A_N(_09234_),
    .B(_08832_),
    .C(_08829_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand3_2 _19571_ (.A(_08829_),
    .B(_09233_),
    .C(_08418_),
    .Y(_09238_));
 sky130_fd_sc_hd__o211a_2 _19572_ (.A1(_08827_),
    .A2(_08828_),
    .B1(_08832_),
    .C1(_09238_),
    .X(_09239_));
 sky130_fd_sc_hd__o211ai_4 _19573_ (.A1(_08827_),
    .A2(_08828_),
    .B1(_08832_),
    .C1(_09238_),
    .Y(_09240_));
 sky130_fd_sc_hd__a31o_2 _19574_ (.A1(_08832_),
    .A2(_08834_),
    .A3(_09238_),
    .B1(_09235_),
    .X(_09241_));
 sky130_fd_sc_hd__o21ai_1 _19575_ (.A1(_09235_),
    .A2(_09239_),
    .B1(_09232_),
    .Y(_09242_));
 sky130_fd_sc_hd__o211ai_1 _19576_ (.A1(_09228_),
    .A2(_09230_),
    .B1(_09237_),
    .C1(_09240_),
    .Y(_09243_));
 sky130_fd_sc_hd__nand4_4 _19577_ (.A(_09229_),
    .B(_09231_),
    .C(_09237_),
    .D(_09240_),
    .Y(_09244_));
 sky130_fd_sc_hd__o22ai_4 _19578_ (.A1(_09228_),
    .A2(_09230_),
    .B1(_09235_),
    .B2(_09239_),
    .Y(_09245_));
 sky130_fd_sc_hd__nand3_1 _19579_ (.A(_09242_),
    .B(_09243_),
    .C(net338),
    .Y(_09246_));
 sky130_fd_sc_hd__and3_1 _19580_ (.A(_08689_),
    .B(_08711_),
    .C(_09227_),
    .X(_09248_));
 sky130_fd_sc_hd__or3_2 _19581_ (.A(_08678_),
    .B(_08700_),
    .C(_09226_),
    .X(_09249_));
 sky130_fd_sc_hd__nand3_2 _19582_ (.A(_09245_),
    .B(net338),
    .C(_09244_),
    .Y(_09250_));
 sky130_fd_sc_hd__a31o_1 _19583_ (.A1(_09245_),
    .A2(net338),
    .A3(_09244_),
    .B1(_09248_),
    .X(_09251_));
 sky130_fd_sc_hd__and3_2 _19584_ (.A(_09251_),
    .B(_09818_),
    .C(_09796_),
    .X(_09252_));
 sky130_fd_sc_hd__a211o_1 _19585_ (.A1(_09249_),
    .A2(_09250_),
    .B1(net351),
    .C1(_09807_),
    .X(_09253_));
 sky130_fd_sc_hd__a311oi_4 _19586_ (.A1(_09245_),
    .A2(net338),
    .A3(_09244_),
    .B1(_09248_),
    .C1(net232),
    .Y(_09254_));
 sky130_fd_sc_hd__nand3_4 _19587_ (.A(_09250_),
    .B(net234),
    .C(_09249_),
    .Y(_09255_));
 sky130_fd_sc_hd__a2bb2oi_1 _19588_ (.A1_N(_06622_),
    .A2_N(_06624_),
    .B1(_09249_),
    .B2(_09250_),
    .Y(_09256_));
 sky130_fd_sc_hd__o211ai_4 _19589_ (.A1(_09227_),
    .A2(net338),
    .B1(net232),
    .C1(_09246_),
    .Y(_09257_));
 sky130_fd_sc_hd__o311a_1 _19590_ (.A1(net286),
    .A2(_06012_),
    .A3(_08431_),
    .B1(_08843_),
    .C1(_08847_),
    .X(_09259_));
 sky130_fd_sc_hd__a31o_1 _19591_ (.A1(_08433_),
    .A2(_08842_),
    .A3(_08845_),
    .B1(_08846_),
    .X(_09260_));
 sky130_fd_sc_hd__a31oi_4 _19592_ (.A1(_08433_),
    .A2(_08842_),
    .A3(_08845_),
    .B1(_08846_),
    .Y(_09261_));
 sky130_fd_sc_hd__a21oi_1 _19593_ (.A1(_09255_),
    .A2(_09257_),
    .B1(_09260_),
    .Y(_09262_));
 sky130_fd_sc_hd__o2bb2ai_2 _19594_ (.A1_N(_09255_),
    .A2_N(_09257_),
    .B1(_09259_),
    .B2(_08844_),
    .Y(_09263_));
 sky130_fd_sc_hd__nor3_1 _19595_ (.A(_09261_),
    .B(_09256_),
    .C(_09254_),
    .Y(_09264_));
 sky130_fd_sc_hd__nand3_2 _19596_ (.A(_09260_),
    .B(_09257_),
    .C(_09255_),
    .Y(_09265_));
 sky130_fd_sc_hd__nand3_1 _19597_ (.A(_09263_),
    .B(_09265_),
    .C(net336),
    .Y(_09266_));
 sky130_fd_sc_hd__o22ai_2 _19598_ (.A1(_09785_),
    .A2(_09807_),
    .B1(_09262_),
    .B2(_09264_),
    .Y(_09267_));
 sky130_fd_sc_hd__a31o_1 _19599_ (.A1(_09263_),
    .A2(_09265_),
    .A3(net336),
    .B1(_09252_),
    .X(_09268_));
 sky130_fd_sc_hd__a2bb2oi_2 _19600_ (.A1_N(_06305_),
    .A2_N(net283),
    .B1(_09253_),
    .B2(_09266_),
    .Y(_09270_));
 sky130_fd_sc_hd__o221ai_4 _19601_ (.A1(_06305_),
    .A2(net283),
    .B1(_09251_),
    .B2(net336),
    .C1(_09267_),
    .Y(_09271_));
 sky130_fd_sc_hd__a31oi_1 _19602_ (.A1(_09263_),
    .A2(_09265_),
    .A3(net336),
    .B1(net251),
    .Y(_09272_));
 sky130_fd_sc_hd__a31o_2 _19603_ (.A1(_09263_),
    .A2(_09265_),
    .A3(net336),
    .B1(net251),
    .X(_09273_));
 sky130_fd_sc_hd__o211a_1 _19604_ (.A1(_06309_),
    .A2(_06312_),
    .B1(_09253_),
    .C1(_09266_),
    .X(_09274_));
 sky130_fd_sc_hd__a311o_1 _19605_ (.A1(_09263_),
    .A2(_09265_),
    .A3(net336),
    .B1(net251),
    .C1(_09252_),
    .X(_09275_));
 sky130_fd_sc_hd__a21oi_1 _19606_ (.A1(_09253_),
    .A2(_09272_),
    .B1(_09270_),
    .Y(_09276_));
 sky130_fd_sc_hd__o32a_1 _19607_ (.A1(net286),
    .A2(_06012_),
    .A3(_08857_),
    .B1(_08862_),
    .B2(_08864_),
    .X(_09277_));
 sky130_fd_sc_hd__o22ai_4 _19608_ (.A1(net254),
    .A2(_08857_),
    .B1(_08862_),
    .B2(_08864_),
    .Y(_09278_));
 sky130_fd_sc_hd__a21oi_1 _19609_ (.A1(_09271_),
    .A2(_09275_),
    .B1(_09278_),
    .Y(_09279_));
 sky130_fd_sc_hd__o21ai_1 _19610_ (.A1(_09270_),
    .A2(_09274_),
    .B1(_09277_),
    .Y(_09281_));
 sky130_fd_sc_hd__o211a_1 _19611_ (.A1(_09273_),
    .A2(_09252_),
    .B1(_09271_),
    .C1(_09278_),
    .X(_09282_));
 sky130_fd_sc_hd__o211ai_1 _19612_ (.A1(_09273_),
    .A2(_09252_),
    .B1(_09271_),
    .C1(_09278_),
    .Y(_09283_));
 sky130_fd_sc_hd__o22ai_2 _19613_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_09279_),
    .B2(_09282_),
    .Y(_09284_));
 sky130_fd_sc_hd__a211o_2 _19614_ (.A1(_09253_),
    .A2(_09266_),
    .B1(_11046_),
    .C1(_11057_),
    .X(_09285_));
 sky130_fd_sc_hd__nand3_2 _19615_ (.A(_09281_),
    .B(_09283_),
    .C(net333),
    .Y(_09286_));
 sky130_fd_sc_hd__a2bb2oi_2 _19616_ (.A1_N(_06009_),
    .A2_N(_06010_),
    .B1(_09285_),
    .B2(_09286_),
    .Y(_09287_));
 sky130_fd_sc_hd__o211ai_2 _19617_ (.A1(_09268_),
    .A2(net333),
    .B1(net253),
    .C1(_09284_),
    .Y(_09288_));
 sky130_fd_sc_hd__o211a_1 _19618_ (.A1(net286),
    .A2(_06012_),
    .B1(_09285_),
    .C1(_09286_),
    .X(_09289_));
 sky130_fd_sc_hd__o211ai_2 _19619_ (.A1(net286),
    .A2(_06012_),
    .B1(_09285_),
    .C1(_09286_),
    .Y(_09290_));
 sky130_fd_sc_hd__o21ai_1 _19620_ (.A1(net261),
    .A2(_08868_),
    .B1(_08883_),
    .Y(_09292_));
 sky130_fd_sc_hd__o22ai_2 _19621_ (.A1(net262),
    .A2(_08869_),
    .B1(_09292_),
    .B2(_08881_),
    .Y(_09293_));
 sky130_fd_sc_hd__a31oi_2 _19622_ (.A1(_08873_),
    .A2(_08882_),
    .A3(_08883_),
    .B1(_08870_),
    .Y(_09294_));
 sky130_fd_sc_hd__nand3_2 _19623_ (.A(_09293_),
    .B(_09290_),
    .C(_09288_),
    .Y(_09295_));
 sky130_fd_sc_hd__o21ai_2 _19624_ (.A1(_09287_),
    .A2(_09289_),
    .B1(_09294_),
    .Y(_09296_));
 sky130_fd_sc_hd__o211a_1 _19625_ (.A1(_09268_),
    .A2(net333),
    .B1(_12703_),
    .C1(_09284_),
    .X(_09297_));
 sky130_fd_sc_hd__a211o_2 _19626_ (.A1(_09285_),
    .A2(_09286_),
    .B1(_12670_),
    .C1(net327),
    .X(_09298_));
 sky130_fd_sc_hd__nand3_2 _19627_ (.A(_09295_),
    .B(_09296_),
    .C(net312),
    .Y(_09299_));
 sky130_fd_sc_hd__a31o_1 _19628_ (.A1(_09295_),
    .A2(_09296_),
    .A3(net312),
    .B1(_09297_),
    .X(_09300_));
 sky130_fd_sc_hd__a31oi_2 _19629_ (.A1(_09295_),
    .A2(_09296_),
    .A3(net312),
    .B1(_09297_),
    .Y(_09301_));
 sky130_fd_sc_hd__and3_4 _19630_ (.A(_09300_),
    .B(_00044_),
    .C(_00022_),
    .X(_09303_));
 sky130_fd_sc_hd__or3_1 _19631_ (.A(net324),
    .B(_00033_),
    .C(_09301_),
    .X(_09304_));
 sky130_fd_sc_hd__nand3_1 _19632_ (.A(_08112_),
    .B(_07739_),
    .C(_08110_),
    .Y(_09305_));
 sky130_fd_sc_hd__a211oi_4 _19633_ (.A1(_08473_),
    .A2(_08493_),
    .B1(_09305_),
    .C1(_08496_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand2_1 _19634_ (.A(_08898_),
    .B(_09306_),
    .Y(_09307_));
 sky130_fd_sc_hd__o211a_1 _19635_ (.A1(_08903_),
    .A2(_08897_),
    .B1(_08899_),
    .C1(_09307_),
    .X(_09308_));
 sky130_fd_sc_hd__o211ai_4 _19636_ (.A1(_08903_),
    .A2(_08897_),
    .B1(_08899_),
    .C1(_09307_),
    .Y(_09309_));
 sky130_fd_sc_hd__nand4_4 _19637_ (.A(_07736_),
    .B(_08898_),
    .C(_08899_),
    .D(_09306_),
    .Y(_09310_));
 sky130_fd_sc_hd__a41o_1 _19638_ (.A1(_07736_),
    .A2(_08898_),
    .A3(_08899_),
    .A4(_09306_),
    .B1(_09308_),
    .X(_09311_));
 sky130_fd_sc_hd__a21oi_4 _19639_ (.A1(_09298_),
    .A2(_09299_),
    .B1(net262),
    .Y(_09312_));
 sky130_fd_sc_hd__o21ai_4 _19640_ (.A1(_05760_),
    .A2(net290),
    .B1(_09300_),
    .Y(_09314_));
 sky130_fd_sc_hd__and3_1 _19641_ (.A(_09299_),
    .B(net262),
    .C(_09298_),
    .X(_09315_));
 sky130_fd_sc_hd__o211ai_4 _19642_ (.A1(_05765_),
    .A2(net289),
    .B1(_09298_),
    .C1(_09299_),
    .Y(_09316_));
 sky130_fd_sc_hd__nor2_1 _19643_ (.A(_09312_),
    .B(_09315_),
    .Y(_09317_));
 sky130_fd_sc_hd__o2bb2ai_4 _19644_ (.A1_N(_09309_),
    .A2_N(_09310_),
    .B1(_09312_),
    .B2(_09315_),
    .Y(_09318_));
 sky130_fd_sc_hd__nand4_4 _19645_ (.A(_09309_),
    .B(_09310_),
    .C(_09314_),
    .D(_09316_),
    .Y(_09319_));
 sky130_fd_sc_hd__nand3_1 _19646_ (.A(_09318_),
    .B(_09319_),
    .C(net309),
    .Y(_09320_));
 sky130_fd_sc_hd__a31oi_4 _19647_ (.A1(_09318_),
    .A2(_09319_),
    .A3(net309),
    .B1(_09303_),
    .Y(_09321_));
 sky130_fd_sc_hd__a31o_1 _19648_ (.A1(_09318_),
    .A2(_09319_),
    .A3(net309),
    .B1(_09303_),
    .X(_09322_));
 sky130_fd_sc_hd__a2bb2o_2 _19649_ (.A1_N(_01919_),
    .A2_N(_01930_),
    .B1(_09304_),
    .B2(_09320_),
    .X(_09323_));
 sky130_fd_sc_hd__inv_2 _19650_ (.A(_09323_),
    .Y(_09325_));
 sky130_fd_sc_hd__a31o_1 _19651_ (.A1(_09318_),
    .A2(_09319_),
    .A3(net309),
    .B1(net291),
    .X(_09326_));
 sky130_fd_sc_hd__a311oi_4 _19652_ (.A1(_09318_),
    .A2(_09319_),
    .A3(net309),
    .B1(net291),
    .C1(_09303_),
    .Y(_09327_));
 sky130_fd_sc_hd__nand3_2 _19653_ (.A(_09320_),
    .B(net267),
    .C(_09304_),
    .Y(_09328_));
 sky130_fd_sc_hd__a2bb2oi_1 _19654_ (.A1_N(_05500_),
    .A2_N(_05503_),
    .B1(_09304_),
    .B2(_09320_),
    .Y(_09329_));
 sky130_fd_sc_hd__o21ai_4 _19655_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_09322_),
    .Y(_09330_));
 sky130_fd_sc_hd__a21o_1 _19656_ (.A1(_08919_),
    .A2(_08916_),
    .B1(_08920_),
    .X(_09331_));
 sky130_fd_sc_hd__a21oi_2 _19657_ (.A1(_08919_),
    .A2(_08916_),
    .B1(_08920_),
    .Y(_09332_));
 sky130_fd_sc_hd__o21a_2 _19658_ (.A1(_09327_),
    .A2(_09329_),
    .B1(_09332_),
    .X(_09333_));
 sky130_fd_sc_hd__o21ai_2 _19659_ (.A1(_09327_),
    .A2(_09329_),
    .B1(_09332_),
    .Y(_09334_));
 sky130_fd_sc_hd__o21ai_2 _19660_ (.A1(net267),
    .A2(_09321_),
    .B1(_09331_),
    .Y(_09336_));
 sky130_fd_sc_hd__o211ai_4 _19661_ (.A1(_09303_),
    .A2(_09326_),
    .B1(_09331_),
    .C1(_09330_),
    .Y(_09337_));
 sky130_fd_sc_hd__o22ai_4 _19662_ (.A1(_01940_),
    .A2(net303),
    .B1(_09327_),
    .B2(_09336_),
    .Y(_09338_));
 sky130_fd_sc_hd__o211ai_2 _19663_ (.A1(_09327_),
    .A2(_09336_),
    .B1(net280),
    .C1(_09334_),
    .Y(_09339_));
 sky130_fd_sc_hd__o22ai_4 _19664_ (.A1(net280),
    .A2(_09321_),
    .B1(_09333_),
    .B2(_09338_),
    .Y(_09340_));
 sky130_fd_sc_hd__o211a_1 _19665_ (.A1(_02137_),
    .A2(_08522_),
    .B1(_08544_),
    .C1(_08935_),
    .X(_09341_));
 sky130_fd_sc_hd__o221a_1 _19666_ (.A1(_02148_),
    .A2(_08521_),
    .B1(net298),
    .B2(_08931_),
    .C1(_08939_),
    .X(_09342_));
 sky130_fd_sc_hd__a31oi_2 _19667_ (.A1(_08523_),
    .A2(_08544_),
    .A3(_08935_),
    .B1(_08936_),
    .Y(_09343_));
 sky130_fd_sc_hd__a31oi_1 _19668_ (.A1(_09334_),
    .A2(_09337_),
    .A3(net279),
    .B1(net293),
    .Y(_09344_));
 sky130_fd_sc_hd__a311oi_4 _19669_ (.A1(_09334_),
    .A2(_09337_),
    .A3(net279),
    .B1(net293),
    .C1(_09325_),
    .Y(_09345_));
 sky130_fd_sc_hd__o221ai_4 _19670_ (.A1(net280),
    .A2(_09321_),
    .B1(_09333_),
    .B2(_09338_),
    .C1(net295),
    .Y(_09347_));
 sky130_fd_sc_hd__a2bb2oi_2 _19671_ (.A1_N(_05242_),
    .A2_N(net317),
    .B1(_09323_),
    .B2(_09339_),
    .Y(_09348_));
 sky130_fd_sc_hd__o21ai_1 _19672_ (.A1(_05242_),
    .A2(net317),
    .B1(_09340_),
    .Y(_09349_));
 sky130_fd_sc_hd__a21oi_1 _19673_ (.A1(_09323_),
    .A2(_09344_),
    .B1(_09348_),
    .Y(_09350_));
 sky130_fd_sc_hd__o211ai_2 _19674_ (.A1(_08936_),
    .A2(_09341_),
    .B1(_09347_),
    .C1(_09349_),
    .Y(_09351_));
 sky130_fd_sc_hd__o22ai_2 _19675_ (.A1(_08934_),
    .A2(_09342_),
    .B1(_09345_),
    .B2(_09348_),
    .Y(_09352_));
 sky130_fd_sc_hd__o211ai_4 _19676_ (.A1(_04008_),
    .A2(net300),
    .B1(_09351_),
    .C1(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__a211o_1 _19677_ (.A1(_09323_),
    .A2(_09339_),
    .B1(_04008_),
    .C1(net300),
    .X(_09354_));
 sky130_fd_sc_hd__nand3_1 _19678_ (.A(_09349_),
    .B(_09343_),
    .C(_09347_),
    .Y(_09355_));
 sky130_fd_sc_hd__o22ai_1 _19679_ (.A1(_08936_),
    .A2(_09341_),
    .B1(_09345_),
    .B2(_09348_),
    .Y(_09356_));
 sky130_fd_sc_hd__nand3_2 _19680_ (.A(_09356_),
    .B(net276),
    .C(_09355_),
    .Y(_09358_));
 sky130_fd_sc_hd__o21ai_4 _19681_ (.A1(net276),
    .A2(_09340_),
    .B1(_09353_),
    .Y(_09359_));
 sky130_fd_sc_hd__o211a_1 _19682_ (.A1(_09340_),
    .A2(net276),
    .B1(net298),
    .C1(_09353_),
    .X(_09360_));
 sky130_fd_sc_hd__o211ai_4 _19683_ (.A1(_09340_),
    .A2(net276),
    .B1(net298),
    .C1(_09353_),
    .Y(_09361_));
 sky130_fd_sc_hd__nand3_4 _19684_ (.A(_09358_),
    .B(net299),
    .C(_09354_),
    .Y(_09362_));
 sky130_fd_sc_hd__inv_2 _19685_ (.A(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__o22a_1 _19686_ (.A1(_08553_),
    .A2(_08954_),
    .B1(_02137_),
    .B2(_08948_),
    .X(_09364_));
 sky130_fd_sc_hd__o21ai_2 _19687_ (.A1(_08952_),
    .A2(_08956_),
    .B1(_08950_),
    .Y(_09365_));
 sky130_fd_sc_hd__a21oi_4 _19688_ (.A1(_09361_),
    .A2(_09362_),
    .B1(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__o2bb2ai_1 _19689_ (.A1_N(_09361_),
    .A2_N(_09362_),
    .B1(_09364_),
    .B2(_08952_),
    .Y(_09367_));
 sky130_fd_sc_hd__nand3_1 _19690_ (.A(_09361_),
    .B(_09362_),
    .C(_09365_),
    .Y(_09369_));
 sky130_fd_sc_hd__a31o_2 _19691_ (.A1(_09361_),
    .A2(_09362_),
    .A3(_09365_),
    .B1(_05234_),
    .X(_09370_));
 sky130_fd_sc_hd__nand3_1 _19692_ (.A(_09367_),
    .B(_09369_),
    .C(net273),
    .Y(_09371_));
 sky130_fd_sc_hd__a211o_1 _19693_ (.A1(_09354_),
    .A2(_09358_),
    .B1(net297),
    .C1(_05232_),
    .X(_09372_));
 sky130_fd_sc_hd__o22ai_4 _19694_ (.A1(net273),
    .A2(_09359_),
    .B1(_09366_),
    .B2(_09370_),
    .Y(_09373_));
 sky130_fd_sc_hd__a22oi_4 _19695_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_09371_),
    .B2(_09372_),
    .Y(_09374_));
 sky130_fd_sc_hd__o21ai_2 _19696_ (.A1(_02049_),
    .A2(_02071_),
    .B1(_09373_),
    .Y(_09375_));
 sky130_fd_sc_hd__o221a_1 _19697_ (.A1(net273),
    .A2(_09359_),
    .B1(_09366_),
    .B2(_09370_),
    .C1(_02137_),
    .X(_09376_));
 sky130_fd_sc_hd__o221ai_4 _19698_ (.A1(net273),
    .A2(_09359_),
    .B1(_09366_),
    .B2(_09370_),
    .C1(_02137_),
    .Y(_09377_));
 sky130_fd_sc_hd__nand4_1 _19699_ (.A(_07795_),
    .B(_07797_),
    .C(_08172_),
    .D(_08175_),
    .Y(_09378_));
 sky130_fd_sc_hd__a21oi_1 _19700_ (.A1(net326),
    .A2(_08566_),
    .B1(_09378_),
    .Y(_09380_));
 sky130_fd_sc_hd__nor3_1 _19701_ (.A(_08572_),
    .B(_09378_),
    .C(_08574_),
    .Y(_09381_));
 sky130_fd_sc_hd__nand3_1 _19702_ (.A(_09380_),
    .B(_08969_),
    .C(_08573_),
    .Y(_09382_));
 sky130_fd_sc_hd__o211ai_4 _19703_ (.A1(_08975_),
    .A2(_08968_),
    .B1(_08971_),
    .C1(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__nand4_4 _19704_ (.A(_08969_),
    .B(_09381_),
    .C(_08971_),
    .D(_07798_),
    .Y(_09384_));
 sky130_fd_sc_hd__nand2_2 _19705_ (.A(_09383_),
    .B(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__nand4_4 _19706_ (.A(_09375_),
    .B(_09377_),
    .C(_09383_),
    .D(_09384_),
    .Y(_09386_));
 sky130_fd_sc_hd__o21ai_4 _19707_ (.A1(_09374_),
    .A2(_09376_),
    .B1(_09385_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand3_2 _19708_ (.A(_09387_),
    .B(net246),
    .C(_09386_),
    .Y(_09388_));
 sky130_fd_sc_hd__and3_4 _19709_ (.A(_05482_),
    .B(_05484_),
    .C(_09373_),
    .X(_09389_));
 sky130_fd_sc_hd__a211o_2 _19710_ (.A1(_09371_),
    .A2(_09372_),
    .B1(_05481_),
    .C1(_05483_),
    .X(_09391_));
 sky130_fd_sc_hd__a31oi_4 _19711_ (.A1(_09387_),
    .A2(net246),
    .A3(_09386_),
    .B1(_09389_),
    .Y(_09392_));
 sky130_fd_sc_hd__a21oi_2 _19712_ (.A1(_09388_),
    .A2(_09391_),
    .B1(net241),
    .Y(_09393_));
 sky130_fd_sc_hd__or3_2 _19713_ (.A(net266),
    .B(_05751_),
    .C(_09392_),
    .X(_09394_));
 sky130_fd_sc_hd__a31o_2 _19714_ (.A1(_09387_),
    .A2(net246),
    .A3(_09386_),
    .B1(net319),
    .X(_09395_));
 sky130_fd_sc_hd__a311oi_4 _19715_ (.A1(_09387_),
    .A2(net246),
    .A3(_09386_),
    .B1(_09389_),
    .C1(net319),
    .Y(_09396_));
 sky130_fd_sc_hd__a22oi_4 _19716_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_09388_),
    .B2(_09391_),
    .Y(_09397_));
 sky130_fd_sc_hd__a22o_1 _19717_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_09388_),
    .B2(_09391_),
    .X(_09398_));
 sky130_fd_sc_hd__o31a_2 _19718_ (.A1(_08585_),
    .A2(_08983_),
    .A3(_08987_),
    .B1(_08986_),
    .X(_09399_));
 sky130_fd_sc_hd__o31a_1 _19719_ (.A1(_08587_),
    .A2(_08982_),
    .A3(_08985_),
    .B1(_08988_),
    .X(_09400_));
 sky130_fd_sc_hd__o21a_1 _19720_ (.A1(_09396_),
    .A2(_09397_),
    .B1(_09400_),
    .X(_09402_));
 sky130_fd_sc_hd__o21ai_4 _19721_ (.A1(_09396_),
    .A2(_09397_),
    .B1(_09400_),
    .Y(_09403_));
 sky130_fd_sc_hd__o21ai_2 _19722_ (.A1(net320),
    .A2(_09392_),
    .B1(_09399_),
    .Y(_09404_));
 sky130_fd_sc_hd__o211ai_4 _19723_ (.A1(_09389_),
    .A2(_09395_),
    .B1(_09399_),
    .C1(_09398_),
    .Y(_09405_));
 sky130_fd_sc_hd__o22ai_2 _19724_ (.A1(net266),
    .A2(_05751_),
    .B1(_09396_),
    .B2(_09404_),
    .Y(_09406_));
 sky130_fd_sc_hd__o211ai_4 _19725_ (.A1(_09396_),
    .A2(_09404_),
    .B1(net241),
    .C1(_09403_),
    .Y(_09407_));
 sky130_fd_sc_hd__o22ai_4 _19726_ (.A1(net241),
    .A2(_09392_),
    .B1(_09402_),
    .B2(_09406_),
    .Y(_09408_));
 sky130_fd_sc_hd__a311o_2 _19727_ (.A1(_09403_),
    .A2(_09405_),
    .A3(net241),
    .B1(net240),
    .C1(_09393_),
    .X(_09409_));
 sky130_fd_sc_hd__o311a_1 _19728_ (.A1(net365),
    .A2(net364),
    .A3(_08597_),
    .B1(_08610_),
    .C1(_09000_),
    .X(_09410_));
 sky130_fd_sc_hd__o22a_1 _19729_ (.A1(_08600_),
    .A2(_08609_),
    .B1(_11309_),
    .B2(_08998_),
    .X(_09411_));
 sky130_fd_sc_hd__o31a_1 _19730_ (.A1(_08600_),
    .A2(_08609_),
    .A3(_08999_),
    .B1(_09002_),
    .X(_09413_));
 sky130_fd_sc_hd__a31o_1 _19731_ (.A1(_08602_),
    .A2(_08610_),
    .A3(_09000_),
    .B1(_09001_),
    .X(_09414_));
 sky130_fd_sc_hd__a31oi_2 _19732_ (.A1(_09403_),
    .A2(_09405_),
    .A3(net241),
    .B1(net326),
    .Y(_09415_));
 sky130_fd_sc_hd__a311oi_4 _19733_ (.A1(_09403_),
    .A2(_09405_),
    .A3(net241),
    .B1(_09393_),
    .C1(net326),
    .Y(_09416_));
 sky130_fd_sc_hd__o221ai_4 _19734_ (.A1(_12867_),
    .A2(_12877_),
    .B1(net241),
    .B2(_09392_),
    .C1(_09407_),
    .Y(_09417_));
 sky130_fd_sc_hd__a2bb2oi_4 _19735_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_09394_),
    .B2(_09407_),
    .Y(_09418_));
 sky130_fd_sc_hd__o21ai_1 _19736_ (.A1(net361),
    .A2(net345),
    .B1(_09408_),
    .Y(_09419_));
 sky130_fd_sc_hd__o211ai_2 _19737_ (.A1(_09001_),
    .A2(_09410_),
    .B1(_09417_),
    .C1(_09419_),
    .Y(_09420_));
 sky130_fd_sc_hd__o22ai_2 _19738_ (.A1(_08999_),
    .A2(_09411_),
    .B1(_09416_),
    .B2(_09418_),
    .Y(_09421_));
 sky130_fd_sc_hd__o211ai_4 _19739_ (.A1(net259),
    .A2(net257),
    .B1(_09420_),
    .C1(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__a211o_4 _19740_ (.A1(_09394_),
    .A2(_09407_),
    .B1(net259),
    .C1(net257),
    .X(_09424_));
 sky130_fd_sc_hd__nand3_1 _19741_ (.A(_09419_),
    .B(_09413_),
    .C(_09417_),
    .Y(_09425_));
 sky130_fd_sc_hd__o22ai_2 _19742_ (.A1(_09001_),
    .A2(_09410_),
    .B1(_09416_),
    .B2(_09418_),
    .Y(_09426_));
 sky130_fd_sc_hd__o211ai_4 _19743_ (.A1(net259),
    .A2(net257),
    .B1(_09425_),
    .C1(_09426_),
    .Y(_09427_));
 sky130_fd_sc_hd__o31a_1 _19744_ (.A1(net259),
    .A2(net257),
    .A3(_09408_),
    .B1(_09422_),
    .X(_09428_));
 sky130_fd_sc_hd__and3_1 _19745_ (.A(_06294_),
    .B(_09424_),
    .C(_09427_),
    .X(_09429_));
 sky130_fd_sc_hd__a2bb2oi_4 _19746_ (.A1_N(_11210_),
    .A2_N(_11232_),
    .B1(_09424_),
    .B2(_09427_),
    .Y(_09430_));
 sky130_fd_sc_hd__o211ai_4 _19747_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_09409_),
    .C1(_09422_),
    .Y(_09431_));
 sky130_fd_sc_hd__o211a_4 _19748_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_09424_),
    .C1(_09427_),
    .X(_09432_));
 sky130_fd_sc_hd__o211ai_4 _19749_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_09424_),
    .C1(_09427_),
    .Y(_09433_));
 sky130_fd_sc_hd__and3_1 _19750_ (.A(_08621_),
    .B(_09016_),
    .C(_09021_),
    .X(_09435_));
 sky130_fd_sc_hd__o21ai_1 _19751_ (.A1(_09018_),
    .A2(_09022_),
    .B1(_09016_),
    .Y(_09436_));
 sky130_fd_sc_hd__a31o_1 _19752_ (.A1(_08621_),
    .A2(_09016_),
    .A3(_09021_),
    .B1(_09018_),
    .X(_09437_));
 sky130_fd_sc_hd__o211ai_4 _19753_ (.A1(_09018_),
    .A2(_09435_),
    .B1(_09433_),
    .C1(_09431_),
    .Y(_09438_));
 sky130_fd_sc_hd__o22ai_4 _19754_ (.A1(_09015_),
    .A2(_09029_),
    .B1(_09430_),
    .B2(_09432_),
    .Y(_09439_));
 sky130_fd_sc_hd__nand3_1 _19755_ (.A(_09439_),
    .B(net212),
    .C(_09438_),
    .Y(_09440_));
 sky130_fd_sc_hd__a22o_1 _19756_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_09424_),
    .B2(_09427_),
    .X(_09441_));
 sky130_fd_sc_hd__o2bb2ai_1 _19757_ (.A1_N(_09431_),
    .A2_N(_09433_),
    .B1(_09435_),
    .B2(_09018_),
    .Y(_09442_));
 sky130_fd_sc_hd__o21ai_1 _19758_ (.A1(_09015_),
    .A2(_09029_),
    .B1(_09431_),
    .Y(_09443_));
 sky130_fd_sc_hd__o221ai_4 _19759_ (.A1(_06291_),
    .A2(_06292_),
    .B1(_09432_),
    .B2(_09443_),
    .C1(_09442_),
    .Y(_09444_));
 sky130_fd_sc_hd__a31oi_2 _19760_ (.A1(_09439_),
    .A2(net212),
    .A3(_09438_),
    .B1(_09429_),
    .Y(_09446_));
 sky130_fd_sc_hd__or3_1 _19761_ (.A(_06608_),
    .B(net237),
    .C(_09446_),
    .X(_09447_));
 sky130_fd_sc_hd__a311oi_4 _19762_ (.A1(_09439_),
    .A2(net212),
    .A3(_09438_),
    .B1(_09429_),
    .C1(_10015_),
    .Y(_09448_));
 sky130_fd_sc_hd__o211ai_4 _19763_ (.A1(net212),
    .A2(_09428_),
    .B1(_09440_),
    .C1(_10025_),
    .Y(_09449_));
 sky130_fd_sc_hd__o211a_1 _19764_ (.A1(net365),
    .A2(net364),
    .B1(_09441_),
    .C1(_09444_),
    .X(_09450_));
 sky130_fd_sc_hd__o211ai_4 _19765_ (.A1(net365),
    .A2(net364),
    .B1(_09441_),
    .C1(_09444_),
    .Y(_09451_));
 sky130_fd_sc_hd__and2_1 _19766_ (.A(_08722_),
    .B(_09033_),
    .X(_09452_));
 sky130_fd_sc_hd__a32oi_4 _19767_ (.A1(_08918_),
    .A2(_09014_),
    .A3(_09025_),
    .B1(_09033_),
    .B2(_08722_),
    .Y(_09453_));
 sky130_fd_sc_hd__a32o_1 _19768_ (.A1(_08918_),
    .A2(_09014_),
    .A3(_09025_),
    .B1(_09033_),
    .B2(_08722_),
    .X(_09454_));
 sky130_fd_sc_hd__o21ai_1 _19769_ (.A1(_09448_),
    .A2(_09450_),
    .B1(_09453_),
    .Y(_09455_));
 sky130_fd_sc_hd__a31oi_2 _19770_ (.A1(_09444_),
    .A2(_10015_),
    .A3(_09441_),
    .B1(_09453_),
    .Y(_09457_));
 sky130_fd_sc_hd__nand2_1 _19771_ (.A(_09457_),
    .B(_09449_),
    .Y(_09458_));
 sky130_fd_sc_hd__nand3_1 _19772_ (.A(_09449_),
    .B(_09451_),
    .C(_09453_),
    .Y(_09459_));
 sky130_fd_sc_hd__o2bb2ai_1 _19773_ (.A1_N(_09449_),
    .A2_N(_09451_),
    .B1(_09452_),
    .B2(_09034_),
    .Y(_09460_));
 sky130_fd_sc_hd__nand3_2 _19774_ (.A(_09460_),
    .B(net211),
    .C(_09459_),
    .Y(_09461_));
 sky130_fd_sc_hd__a311o_2 _19775_ (.A1(_09439_),
    .A2(net212),
    .A3(_09438_),
    .B1(net211),
    .C1(_09429_),
    .X(_09462_));
 sky130_fd_sc_hd__nand3_2 _19776_ (.A(_09455_),
    .B(_09458_),
    .C(net211),
    .Y(_09463_));
 sky130_fd_sc_hd__o211ai_4 _19777_ (.A1(_08863_),
    .A2(_08885_),
    .B1(_09462_),
    .C1(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__o311a_1 _19778_ (.A1(_06608_),
    .A2(net237),
    .A3(_09446_),
    .B1(_09461_),
    .C1(_08918_),
    .X(_09465_));
 sky130_fd_sc_hd__o211ai_2 _19779_ (.A1(_08819_),
    .A2(_08841_),
    .B1(_09447_),
    .C1(_09461_),
    .Y(_09466_));
 sky130_fd_sc_hd__nand3_4 _19780_ (.A(_09132_),
    .B(_09464_),
    .C(_09466_),
    .Y(_09468_));
 sky130_fd_sc_hd__a21o_2 _19781_ (.A1(_09464_),
    .A2(_09466_),
    .B1(_09132_),
    .X(_09469_));
 sky130_fd_sc_hd__nand3_1 _19782_ (.A(_09469_),
    .B(net208),
    .C(_09468_),
    .Y(_09470_));
 sky130_fd_sc_hd__o311a_2 _19783_ (.A1(_06608_),
    .A2(net237),
    .A3(_09446_),
    .B1(_09461_),
    .C1(_06904_),
    .X(_09471_));
 sky130_fd_sc_hd__a211o_1 _19784_ (.A1(_09462_),
    .A2(_09463_),
    .B1(net230),
    .C1(_06901_),
    .X(_09472_));
 sky130_fd_sc_hd__a31oi_4 _19785_ (.A1(_09469_),
    .A2(net208),
    .A3(_09468_),
    .B1(_09471_),
    .Y(_09473_));
 sky130_fd_sc_hd__a311o_1 _19786_ (.A1(_09469_),
    .A2(net208),
    .A3(_09468_),
    .B1(_09471_),
    .C1(net185),
    .X(_09474_));
 sky130_fd_sc_hd__o32a_1 _19787_ (.A1(_06989_),
    .A2(net375),
    .A3(_09057_),
    .B1(_09062_),
    .B2(_08660_),
    .X(_09475_));
 sky130_fd_sc_hd__o211a_1 _19788_ (.A1(_08665_),
    .A2(_08662_),
    .B1(_08661_),
    .C1(_09065_),
    .X(_09476_));
 sky130_fd_sc_hd__a32o_1 _19789_ (.A1(_09057_),
    .A2(_06978_),
    .A3(_06956_),
    .B1(_09063_),
    .B2(_09067_),
    .X(_09477_));
 sky130_fd_sc_hd__a311oi_4 _19790_ (.A1(_09469_),
    .A2(net208),
    .A3(_09468_),
    .B1(_09471_),
    .C1(_07899_),
    .Y(_09479_));
 sky130_fd_sc_hd__nand3_1 _19791_ (.A(_09470_),
    .B(_09472_),
    .C(_07888_),
    .Y(_09480_));
 sky130_fd_sc_hd__a21oi_2 _19792_ (.A1(_09470_),
    .A2(_09472_),
    .B1(_07888_),
    .Y(_09481_));
 sky130_fd_sc_hd__a22o_1 _19793_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_09470_),
    .B2(_09472_),
    .X(_09482_));
 sky130_fd_sc_hd__o211ai_1 _19794_ (.A1(_09064_),
    .A2(_09475_),
    .B1(_09480_),
    .C1(_09482_),
    .Y(_09483_));
 sky130_fd_sc_hd__o22ai_1 _19795_ (.A1(_09066_),
    .A2(_09476_),
    .B1(_09479_),
    .B2(_09481_),
    .Y(_09484_));
 sky130_fd_sc_hd__nand3_1 _19796_ (.A(net185),
    .B(_09483_),
    .C(_09484_),
    .Y(_09485_));
 sky130_fd_sc_hd__or3_1 _19797_ (.A(_07227_),
    .B(net203),
    .C(_09473_),
    .X(_09486_));
 sky130_fd_sc_hd__o21ai_1 _19798_ (.A1(_09066_),
    .A2(_09476_),
    .B1(_09480_),
    .Y(_09487_));
 sky130_fd_sc_hd__o22ai_2 _19799_ (.A1(_09064_),
    .A2(_09475_),
    .B1(_09479_),
    .B2(_09481_),
    .Y(_09488_));
 sky130_fd_sc_hd__o211ai_4 _19800_ (.A1(_09487_),
    .A2(_09481_),
    .B1(net185),
    .C1(_09488_),
    .Y(_09490_));
 sky130_fd_sc_hd__o21ai_1 _19801_ (.A1(net185),
    .A2(_09473_),
    .B1(_09490_),
    .Y(_09491_));
 sky130_fd_sc_hd__a211o_2 _19802_ (.A1(_09486_),
    .A2(_09490_),
    .B1(_07544_),
    .C1(net184),
    .X(_09492_));
 sky130_fd_sc_hd__o21ai_1 _19803_ (.A1(_09080_),
    .A2(_09078_),
    .B1(_09076_),
    .Y(_09493_));
 sky130_fd_sc_hd__o221a_1 _19804_ (.A1(_06989_),
    .A2(net375),
    .B1(net185),
    .B2(_09473_),
    .C1(_09490_),
    .X(_09494_));
 sky130_fd_sc_hd__o221ai_4 _19805_ (.A1(_06989_),
    .A2(net375),
    .B1(net185),
    .B2(_09473_),
    .C1(_09490_),
    .Y(_09495_));
 sky130_fd_sc_hd__a2bb2oi_1 _19806_ (.A1_N(_06945_),
    .A2_N(_06967_),
    .B1(_09486_),
    .B2(_09490_),
    .Y(_09496_));
 sky130_fd_sc_hd__o211ai_4 _19807_ (.A1(_06945_),
    .A2(_06967_),
    .B1(_09474_),
    .C1(_09485_),
    .Y(_09497_));
 sky130_fd_sc_hd__a32o_1 _19808_ (.A1(_07044_),
    .A2(_09474_),
    .A3(_09485_),
    .B1(_09076_),
    .B2(_09086_),
    .X(_09498_));
 sky130_fd_sc_hd__o211a_1 _19809_ (.A1(_09075_),
    .A2(_09085_),
    .B1(_09495_),
    .C1(_09497_),
    .X(_09499_));
 sky130_fd_sc_hd__a21oi_1 _19810_ (.A1(_09495_),
    .A2(_09497_),
    .B1(_09493_),
    .Y(_09501_));
 sky130_fd_sc_hd__a21o_1 _19811_ (.A1(_09495_),
    .A2(_09497_),
    .B1(_09493_),
    .X(_09502_));
 sky130_fd_sc_hd__o221ai_4 _19812_ (.A1(_07544_),
    .A2(net184),
    .B1(_09494_),
    .B2(_09498_),
    .C1(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__o22ai_2 _19813_ (.A1(_07544_),
    .A2(net184),
    .B1(_09499_),
    .B2(_09501_),
    .Y(_09504_));
 sky130_fd_sc_hd__o21ai_2 _19814_ (.A1(net163),
    .A2(_09491_),
    .B1(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__or3_2 _19815_ (.A(_07912_),
    .B(_07914_),
    .C(_09505_),
    .X(_09506_));
 sky130_fd_sc_hd__a2bb2oi_4 _19816_ (.A1_N(net394),
    .A2_N(_06267_),
    .B1(_09492_),
    .B2(_09503_),
    .Y(_09507_));
 sky130_fd_sc_hd__o211ai_1 _19817_ (.A1(net163),
    .A2(_09491_),
    .B1(_09504_),
    .C1(_06343_),
    .Y(_09508_));
 sky130_fd_sc_hd__o311a_1 _19818_ (.A1(_07550_),
    .A2(_09499_),
    .A3(_09501_),
    .B1(_09492_),
    .C1(_06332_),
    .X(_09509_));
 sky130_fd_sc_hd__o211ai_1 _19819_ (.A1(net381),
    .A2(_06310_),
    .B1(_09492_),
    .C1(_09503_),
    .Y(_09510_));
 sky130_fd_sc_hd__a31o_2 _19820_ (.A1(_09074_),
    .A2(_09087_),
    .A3(_09095_),
    .B1(_09092_),
    .X(_09512_));
 sky130_fd_sc_hd__a21o_1 _19821_ (.A1(_09508_),
    .A2(_09510_),
    .B1(_09512_),
    .X(_09513_));
 sky130_fd_sc_hd__nand3_1 _19822_ (.A(_09508_),
    .B(_09510_),
    .C(_09512_),
    .Y(_09514_));
 sky130_fd_sc_hd__o21ai_1 _19823_ (.A1(_09507_),
    .A2(_09509_),
    .B1(_09512_),
    .Y(_09515_));
 sky130_fd_sc_hd__a31oi_2 _19824_ (.A1(_09503_),
    .A2(_06332_),
    .A3(_09492_),
    .B1(_09512_),
    .Y(_09516_));
 sky130_fd_sc_hd__a31o_1 _19825_ (.A1(_09503_),
    .A2(_06332_),
    .A3(_09492_),
    .B1(_09512_),
    .X(_09517_));
 sky130_fd_sc_hd__o221ai_4 _19826_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_09507_),
    .B2(_09517_),
    .C1(_09515_),
    .Y(_09518_));
 sky130_fd_sc_hd__nand3_1 _19827_ (.A(_09513_),
    .B(_09514_),
    .C(net160),
    .Y(_09519_));
 sky130_fd_sc_hd__o21ai_1 _19828_ (.A1(_07909_),
    .A2(_07911_),
    .B1(_09505_),
    .Y(_09520_));
 sky130_fd_sc_hd__o311ai_4 _19829_ (.A1(_09096_),
    .A2(_09089_),
    .A3(_09088_),
    .B1(_09102_),
    .C1(_09098_),
    .Y(_09521_));
 sky130_fd_sc_hd__and3_2 _19830_ (.A(_09521_),
    .B(_05851_),
    .C(_09103_),
    .X(_09523_));
 sky130_fd_sc_hd__a21oi_2 _19831_ (.A1(_09103_),
    .A2(_09521_),
    .B1(_05851_),
    .Y(_09524_));
 sky130_fd_sc_hd__a22o_1 _19832_ (.A1(net395),
    .A2(_05796_),
    .B1(_09103_),
    .B2(_09521_),
    .X(_09525_));
 sky130_fd_sc_hd__nor3_1 _19833_ (.A(_09524_),
    .B(_08301_),
    .C(_09523_),
    .Y(_09526_));
 sky130_fd_sc_hd__o311a_1 _19834_ (.A1(_08301_),
    .A2(_09523_),
    .A3(_09524_),
    .B1(_09506_),
    .C1(_09518_),
    .X(_09527_));
 sky130_fd_sc_hd__o311ai_4 _19835_ (.A1(_08301_),
    .A2(_09523_),
    .A3(_09524_),
    .B1(_09506_),
    .C1(_09518_),
    .Y(_09528_));
 sky130_fd_sc_hd__and3_1 _19836_ (.A(_09519_),
    .B(_09526_),
    .C(_09520_),
    .X(_09529_));
 sky130_fd_sc_hd__nand3_2 _19837_ (.A(_09519_),
    .B(_09526_),
    .C(_09520_),
    .Y(_09530_));
 sky130_fd_sc_hd__o32ai_4 _19838_ (.A1(_05250_),
    .A2(_09107_),
    .A3(_09109_),
    .B1(_08702_),
    .B2(_09113_),
    .Y(_09531_));
 sky130_fd_sc_hd__o21ai_4 _19839_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__o311a_1 _19840_ (.A1(_05447_),
    .A2(_05469_),
    .A3(_09531_),
    .B1(_08714_),
    .C1(_09532_),
    .X(_09534_));
 sky130_fd_sc_hd__o311ai_4 _19841_ (.A1(_05447_),
    .A2(_05469_),
    .A3(_09531_),
    .B1(_09532_),
    .C1(_08714_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand3_4 _19842_ (.A(_09534_),
    .B(_09530_),
    .C(_09528_),
    .Y(_09536_));
 sky130_fd_sc_hd__o21ai_4 _19843_ (.A1(_09527_),
    .A2(_09529_),
    .B1(_09535_),
    .Y(_09537_));
 sky130_fd_sc_hd__o31ai_1 _19844_ (.A1(_09527_),
    .A2(_09529_),
    .A3(_09535_),
    .B1(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__nand4_1 _19845_ (.A(_05207_),
    .B(_05229_),
    .C(_09536_),
    .D(_09537_),
    .Y(_09539_));
 sky130_fd_sc_hd__a21oi_2 _19846_ (.A1(_09536_),
    .A2(_09537_),
    .B1(_05239_),
    .Y(_09540_));
 sky130_fd_sc_hd__o21ai_2 _19847_ (.A1(net407),
    .A2(_05218_),
    .B1(_09538_),
    .Y(_09541_));
 sky130_fd_sc_hd__nand2_1 _19848_ (.A(_09539_),
    .B(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__a31oi_4 _19849_ (.A1(_09536_),
    .A2(_09537_),
    .A3(_05239_),
    .B1(_09128_),
    .Y(_09543_));
 sky130_fd_sc_hd__a31o_1 _19850_ (.A1(_09536_),
    .A2(_09537_),
    .A3(_05239_),
    .B1(_09128_),
    .X(_09545_));
 sky130_fd_sc_hd__a22oi_1 _19851_ (.A1(_09541_),
    .A2(_09543_),
    .B1(_09542_),
    .B2(_09128_),
    .Y(_09546_));
 sky130_fd_sc_hd__a21oi_1 _19852_ (.A1(_09536_),
    .A2(_09537_),
    .B1(_09125_),
    .Y(_09547_));
 sky130_fd_sc_hd__a21oi_1 _19853_ (.A1(_09546_),
    .A2(_09125_),
    .B1(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__a211o_1 _19854_ (.A1(_09546_),
    .A2(_09125_),
    .B1(_03289_),
    .C1(_09547_),
    .X(_09549_));
 sky130_fd_sc_hd__or2_1 _19855_ (.A(net1),
    .B(_09548_),
    .X(_09550_));
 sky130_fd_sc_hd__nor2_8 _19856_ (.A(net50),
    .B(_09118_),
    .Y(_09551_));
 sky130_fd_sc_hd__or4_4 _19857_ (.A(net48),
    .B(net49),
    .C(net50),
    .D(_08292_),
    .X(_09552_));
 sky130_fd_sc_hd__and3b_4 _19858_ (.A_N(net51),
    .B(_09552_),
    .C(net409),
    .X(_09553_));
 sky130_fd_sc_hd__or3b_2 _19859_ (.A(net51),
    .B(_09551_),
    .C_N(net409),
    .X(_09554_));
 sky130_fd_sc_hd__a21boi_4 _19860_ (.A1(_09552_),
    .A2(net409),
    .B1_N(net51),
    .Y(_09556_));
 sky130_fd_sc_hd__a21bo_1 _19861_ (.A1(_09552_),
    .A2(net409),
    .B1_N(net51),
    .X(_09557_));
 sky130_fd_sc_hd__nand2_8 _19862_ (.A(net409),
    .B(net51),
    .Y(_09558_));
 sky130_fd_sc_hd__o311a_4 _19863_ (.A1(net49),
    .A2(net50),
    .A3(_08704_),
    .B1(net51),
    .C1(net409),
    .X(_09559_));
 sky130_fd_sc_hd__a21oi_4 _19864_ (.A1(_09552_),
    .A2(net409),
    .B1(net51),
    .Y(_09560_));
 sky130_fd_sc_hd__a21o_4 _19865_ (.A1(_09552_),
    .A2(net409),
    .B1(net51),
    .X(_09561_));
 sky130_fd_sc_hd__o21ai_4 _19866_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__o21a_4 _19867_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .X(_09563_));
 sky130_fd_sc_hd__and3_1 _19868_ (.A(_09549_),
    .B(_09550_),
    .C(net143),
    .X(_09564_));
 sky130_fd_sc_hd__a21oi_1 _19869_ (.A1(_09548_),
    .A2(_09562_),
    .B1(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__o21ai_1 _19870_ (.A1(_05051_),
    .A2(_09130_),
    .B1(_09565_),
    .Y(_09567_));
 sky130_fd_sc_hd__or3_1 _19871_ (.A(_05051_),
    .B(_09130_),
    .C(_09565_),
    .X(_09568_));
 sky130_fd_sc_hd__and2_1 _19872_ (.A(_09567_),
    .B(_09568_),
    .X(net83));
 sky130_fd_sc_hd__o2bb2a_1 _19873_ (.A1_N(_09130_),
    .A2_N(_09565_),
    .B1(_04832_),
    .B2(_04942_),
    .X(_09569_));
 sky130_fd_sc_hd__o21ai_4 _19874_ (.A1(net51),
    .A2(_09552_),
    .B1(net409),
    .Y(_09570_));
 sky130_fd_sc_hd__nor2_8 _19875_ (.A(net52),
    .B(_09570_),
    .Y(_09571_));
 sky130_fd_sc_hd__clkinv_4 _19876_ (.A(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__and2_4 _19877_ (.A(_09570_),
    .B(net52),
    .X(_09573_));
 sky130_fd_sc_hd__clkinv_4 _19878_ (.A(_09573_),
    .Y(_09574_));
 sky130_fd_sc_hd__nand2b_4 _19879_ (.A_N(net52),
    .B(_09570_),
    .Y(_09575_));
 sky130_fd_sc_hd__o211ai_4 _19880_ (.A1(net51),
    .A2(_09552_),
    .B1(net52),
    .C1(net409),
    .Y(_09577_));
 sky130_fd_sc_hd__nand2_8 _19881_ (.A(_09575_),
    .B(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__or2_4 _19882_ (.A(_09571_),
    .B(_09573_),
    .X(_09579_));
 sky130_fd_sc_hd__o311a_1 _19883_ (.A1(net381),
    .A2(_06310_),
    .A3(_09073_),
    .B1(_09086_),
    .C1(_09497_),
    .X(_09580_));
 sky130_fd_sc_hd__a32o_1 _19884_ (.A1(_09490_),
    .A2(_07033_),
    .A3(_09486_),
    .B1(_09076_),
    .B2(_09086_),
    .X(_09581_));
 sky130_fd_sc_hd__a21o_1 _19885_ (.A1(_09493_),
    .A2(_09495_),
    .B1(_09496_),
    .X(_09582_));
 sky130_fd_sc_hd__a31oi_2 _19886_ (.A1(_09463_),
    .A2(_08907_),
    .A3(_09462_),
    .B1(_09131_),
    .Y(_09583_));
 sky130_fd_sc_hd__a21oi_1 _19887_ (.A1(_09132_),
    .A2(_09464_),
    .B1(_09465_),
    .Y(_09584_));
 sky130_fd_sc_hd__a32o_1 _19888_ (.A1(_08918_),
    .A2(_09447_),
    .A3(_09461_),
    .B1(_09464_),
    .B2(_09132_),
    .X(_09585_));
 sky130_fd_sc_hd__or4_4 _19889_ (.A(net17),
    .B(net18),
    .C(net19),
    .D(_08306_),
    .X(_09586_));
 sky130_fd_sc_hd__and3b_4 _19890_ (.A_N(net20),
    .B(_09586_),
    .C(net410),
    .X(_09588_));
 sky130_fd_sc_hd__or3b_4 _19891_ (.A(_03399_),
    .B(net20),
    .C_N(_09586_),
    .X(_09589_));
 sky130_fd_sc_hd__a21boi_4 _19892_ (.A1(_09586_),
    .A2(net410),
    .B1_N(net20),
    .Y(_09590_));
 sky130_fd_sc_hd__a21bo_4 _19893_ (.A1(_09586_),
    .A2(net410),
    .B1_N(net20),
    .X(_09591_));
 sky130_fd_sc_hd__a21oi_4 _19894_ (.A1(_09586_),
    .A2(net410),
    .B1(net20),
    .Y(_09592_));
 sky130_fd_sc_hd__o311a_4 _19895_ (.A1(net18),
    .A2(net19),
    .A3(_08723_),
    .B1(net20),
    .C1(net410),
    .X(_09593_));
 sky130_fd_sc_hd__nor2_8 _19896_ (.A(net189),
    .B(net186),
    .Y(_09594_));
 sky130_fd_sc_hd__nor2_8 _19897_ (.A(_09592_),
    .B(_09593_),
    .Y(_09595_));
 sky130_fd_sc_hd__o221a_1 _19898_ (.A1(_05130_),
    .A2(_05152_),
    .B1(_09588_),
    .B2(_09590_),
    .C1(net33),
    .X(_09596_));
 sky130_fd_sc_hd__a211o_1 _19899_ (.A1(_09595_),
    .A2(net33),
    .B1(_09134_),
    .C1(_09135_),
    .X(_09597_));
 sky130_fd_sc_hd__o21ai_2 _19900_ (.A1(_09142_),
    .A2(net172),
    .B1(_09597_),
    .Y(_09599_));
 sky130_fd_sc_hd__inv_2 _19901_ (.A(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__o22ai_4 _19902_ (.A1(_08733_),
    .A2(net174),
    .B1(_09145_),
    .B2(_09143_),
    .Y(_09601_));
 sky130_fd_sc_hd__nand2_1 _19903_ (.A(_09601_),
    .B(_09600_),
    .Y(_09602_));
 sky130_fd_sc_hd__o221ai_4 _19904_ (.A1(_08733_),
    .A2(net174),
    .B1(_09145_),
    .B2(_09143_),
    .C1(_09599_),
    .Y(_09603_));
 sky130_fd_sc_hd__o32a_1 _19905_ (.A1(_09593_),
    .A2(_03178_),
    .A3(_09592_),
    .B1(_05130_),
    .B2(_05152_),
    .X(_09604_));
 sky130_fd_sc_hd__a21oi_1 _19906_ (.A1(_09602_),
    .A2(_09603_),
    .B1(_05185_),
    .Y(_09605_));
 sky130_fd_sc_hd__a31oi_4 _19907_ (.A1(_09602_),
    .A2(_09603_),
    .A3(net405),
    .B1(_09596_),
    .Y(_09606_));
 sky130_fd_sc_hd__nor2_2 _19908_ (.A(_05403_),
    .B(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__a311o_1 _19909_ (.A1(_09602_),
    .A2(_09603_),
    .A3(net405),
    .B1(net175),
    .C1(_09596_),
    .X(_09608_));
 sky130_fd_sc_hd__a21o_2 _19910_ (.A1(_08725_),
    .A2(_08727_),
    .B1(_09606_),
    .X(_09610_));
 sky130_fd_sc_hd__o41a_2 _19911_ (.A1(_08728_),
    .A2(net195),
    .A3(_09604_),
    .A4(_09605_),
    .B1(_09608_),
    .X(_09611_));
 sky130_fd_sc_hd__nand2_2 _19912_ (.A(_09608_),
    .B(_09610_),
    .Y(_09612_));
 sky130_fd_sc_hd__o22ai_2 _19913_ (.A1(net199),
    .A2(_09153_),
    .B1(_09162_),
    .B2(_09165_),
    .Y(_09613_));
 sky130_fd_sc_hd__o21a_1 _19914_ (.A1(net198),
    .A2(_09152_),
    .B1(_09163_),
    .X(_09614_));
 sky130_fd_sc_hd__o21ai_1 _19915_ (.A1(net198),
    .A2(_09152_),
    .B1(_09163_),
    .Y(_09615_));
 sky130_fd_sc_hd__a21oi_2 _19916_ (.A1(_09166_),
    .A2(_09614_),
    .B1(_09156_),
    .Y(_09616_));
 sky130_fd_sc_hd__o211a_1 _19917_ (.A1(net198),
    .A2(_09152_),
    .B1(_09611_),
    .C1(_09613_),
    .X(_09617_));
 sky130_fd_sc_hd__o211ai_4 _19918_ (.A1(net198),
    .A2(_09152_),
    .B1(_09611_),
    .C1(_09613_),
    .Y(_09618_));
 sky130_fd_sc_hd__o211ai_2 _19919_ (.A1(_09615_),
    .A2(_09165_),
    .B1(_09157_),
    .C1(_09612_),
    .Y(_09619_));
 sky130_fd_sc_hd__o21ai_2 _19920_ (.A1(_05348_),
    .A2(net401),
    .B1(_09619_),
    .Y(_09621_));
 sky130_fd_sc_hd__o22ai_4 _19921_ (.A1(_05403_),
    .A2(_09606_),
    .B1(_09621_),
    .B2(_09617_),
    .Y(_09622_));
 sky130_fd_sc_hd__inv_2 _19922_ (.A(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__o21a_1 _19923_ (.A1(_08307_),
    .A2(_08309_),
    .B1(_09622_),
    .X(_09624_));
 sky130_fd_sc_hd__o21ai_4 _19924_ (.A1(_08307_),
    .A2(_08309_),
    .B1(_09622_),
    .Y(_09625_));
 sky130_fd_sc_hd__a31o_1 _19925_ (.A1(_05403_),
    .A2(_09618_),
    .A3(_09619_),
    .B1(net198),
    .X(_09626_));
 sky130_fd_sc_hd__nor2_1 _19926_ (.A(net198),
    .B(_09622_),
    .Y(_09627_));
 sky130_fd_sc_hd__a311o_1 _19927_ (.A1(_05403_),
    .A2(_09618_),
    .A3(_09619_),
    .B1(net198),
    .C1(_09607_),
    .X(_09628_));
 sky130_fd_sc_hd__o21a_1 _19928_ (.A1(_09607_),
    .A2(_09626_),
    .B1(_09625_),
    .X(_09629_));
 sky130_fd_sc_hd__o21ai_1 _19929_ (.A1(_09607_),
    .A2(_09626_),
    .B1(_09625_),
    .Y(_09630_));
 sky130_fd_sc_hd__o2111ai_2 _19930_ (.A1(_08351_),
    .A2(_08329_),
    .B1(_07970_),
    .C1(_07968_),
    .D1(_08350_),
    .Y(_09632_));
 sky130_fd_sc_hd__nor3b_2 _19931_ (.A(_08767_),
    .B(_09632_),
    .C_N(_08769_),
    .Y(_09633_));
 sky130_fd_sc_hd__nand4_1 _19932_ (.A(_08768_),
    .B(_08769_),
    .C(_07971_),
    .D(_08352_),
    .Y(_09634_));
 sky130_fd_sc_hd__a21oi_1 _19933_ (.A1(_09633_),
    .A2(_09182_),
    .B1(_09177_),
    .Y(_09635_));
 sky130_fd_sc_hd__o21ai_1 _19934_ (.A1(_09634_),
    .A2(_09180_),
    .B1(_09178_),
    .Y(_09636_));
 sky130_fd_sc_hd__a21oi_4 _19935_ (.A1(_09186_),
    .A2(_09183_),
    .B1(_09636_),
    .Y(_09637_));
 sky130_fd_sc_hd__o21ai_2 _19936_ (.A1(_09184_),
    .A2(_09185_),
    .B1(_09635_),
    .Y(_09638_));
 sky130_fd_sc_hd__and3_1 _19937_ (.A(_09183_),
    .B(_09633_),
    .C(_07982_),
    .X(_09639_));
 sky130_fd_sc_hd__nand4_4 _19938_ (.A(_09178_),
    .B(_09633_),
    .C(_09182_),
    .D(_07982_),
    .Y(_09640_));
 sky130_fd_sc_hd__o31a_1 _19939_ (.A1(_07981_),
    .A2(_09184_),
    .A3(_09634_),
    .B1(_09638_),
    .X(_09641_));
 sky130_fd_sc_hd__o211ai_4 _19940_ (.A1(_09626_),
    .A2(_09607_),
    .B1(_09625_),
    .C1(_09640_),
    .Y(_09643_));
 sky130_fd_sc_hd__a21oi_1 _19941_ (.A1(_09187_),
    .A2(_09635_),
    .B1(_09643_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand3_4 _19942_ (.A(_09638_),
    .B(_09640_),
    .C(_09629_),
    .Y(_09645_));
 sky130_fd_sc_hd__a22oi_2 _19943_ (.A1(_09625_),
    .A2(_09628_),
    .B1(_09638_),
    .B2(_09640_),
    .Y(_09646_));
 sky130_fd_sc_hd__o22ai_4 _19944_ (.A1(_09624_),
    .A2(_09627_),
    .B1(_09637_),
    .B2(_09639_),
    .Y(_09647_));
 sky130_fd_sc_hd__nand3_2 _19945_ (.A(_09647_),
    .B(net358),
    .C(_09645_),
    .Y(_09648_));
 sky130_fd_sc_hd__o21ai_4 _19946_ (.A1(_05654_),
    .A2(_05665_),
    .B1(_09622_),
    .Y(_09649_));
 sky130_fd_sc_hd__inv_2 _19947_ (.A(_09649_),
    .Y(_09650_));
 sky130_fd_sc_hd__o221a_1 _19948_ (.A1(_05403_),
    .A2(_09606_),
    .B1(_09621_),
    .B2(_09617_),
    .C1(_05731_),
    .X(_09651_));
 sky130_fd_sc_hd__a2bb2oi_1 _19949_ (.A1_N(_05676_),
    .A2_N(_05698_),
    .B1(_09645_),
    .B2(_09647_),
    .Y(_09652_));
 sky130_fd_sc_hd__o22ai_2 _19950_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_09644_),
    .B2(_09646_),
    .Y(_09654_));
 sky130_fd_sc_hd__a31oi_4 _19951_ (.A1(_09647_),
    .A2(net358),
    .A3(_09645_),
    .B1(_09650_),
    .Y(_09655_));
 sky130_fd_sc_hd__or4_4 _19952_ (.A(net379),
    .B(net378),
    .C(_09651_),
    .D(_09652_),
    .X(_09656_));
 sky130_fd_sc_hd__o221ai_4 _19953_ (.A1(_07564_),
    .A2(_09191_),
    .B1(_08789_),
    .B2(_08790_),
    .C1(_08785_),
    .Y(_09657_));
 sky130_fd_sc_hd__a31oi_1 _19954_ (.A1(_08785_),
    .A2(_08793_),
    .A3(_09194_),
    .B1(_09195_),
    .Y(_09658_));
 sky130_fd_sc_hd__a311oi_4 _19955_ (.A1(_09647_),
    .A2(net358),
    .A3(_09645_),
    .B1(_09650_),
    .C1(_07936_),
    .Y(_09659_));
 sky130_fd_sc_hd__nand3_4 _19956_ (.A(_09648_),
    .B(_09649_),
    .C(_07935_),
    .Y(_09660_));
 sky130_fd_sc_hd__a22oi_4 _19957_ (.A1(_07929_),
    .A2(_07932_),
    .B1(_09648_),
    .B2(_09649_),
    .Y(_09661_));
 sky130_fd_sc_hd__o211ai_4 _19958_ (.A1(_09622_),
    .A2(net358),
    .B1(_07936_),
    .C1(_09654_),
    .Y(_09662_));
 sky130_fd_sc_hd__nand4_4 _19959_ (.A(_09196_),
    .B(_09657_),
    .C(_09660_),
    .D(_09662_),
    .Y(_09663_));
 sky130_fd_sc_hd__o2bb2ai_4 _19960_ (.A1_N(_09196_),
    .A2_N(_09657_),
    .B1(_09659_),
    .B2(_09661_),
    .Y(_09665_));
 sky130_fd_sc_hd__o211ai_4 _19961_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_09663_),
    .C1(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__o311a_2 _19962_ (.A1(_05731_),
    .A2(_09644_),
    .A3(_09646_),
    .B1(_09649_),
    .C1(_06848_),
    .X(_09667_));
 sky130_fd_sc_hd__a2bb2oi_2 _19963_ (.A1_N(_06793_),
    .A2_N(_06815_),
    .B1(_09663_),
    .B2(_09665_),
    .Y(_09668_));
 sky130_fd_sc_hd__o21ai_1 _19964_ (.A1(net357),
    .A2(_09655_),
    .B1(_09666_),
    .Y(_09669_));
 sky130_fd_sc_hd__a21oi_2 _19965_ (.A1(_09656_),
    .A2(_09666_),
    .B1(net355),
    .Y(_09670_));
 sky130_fd_sc_hd__inv_2 _19966_ (.A(_09670_),
    .Y(_09671_));
 sky130_fd_sc_hd__a2bb2oi_4 _19967_ (.A1_N(_07555_),
    .A2_N(net218),
    .B1(_09656_),
    .B2(_09666_),
    .Y(_09672_));
 sky130_fd_sc_hd__a22o_2 _19968_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_09656_),
    .B2(_09666_),
    .X(_09673_));
 sky130_fd_sc_hd__a31oi_2 _19969_ (.A1(_09663_),
    .A2(_09665_),
    .A3(net357),
    .B1(net202),
    .Y(_09674_));
 sky130_fd_sc_hd__and3_1 _19970_ (.A(_09666_),
    .B(_07564_),
    .C(_09656_),
    .X(_09676_));
 sky130_fd_sc_hd__o211ai_2 _19971_ (.A1(net357),
    .A2(_09655_),
    .B1(_07564_),
    .C1(_09666_),
    .Y(_09677_));
 sky130_fd_sc_hd__a21oi_4 _19972_ (.A1(_09656_),
    .A2(_09674_),
    .B1(_09672_),
    .Y(_09678_));
 sky130_fd_sc_hd__o41ai_4 _19973_ (.A1(_07560_),
    .A2(_07562_),
    .A3(_09667_),
    .A4(_09668_),
    .B1(_09677_),
    .Y(_09679_));
 sky130_fd_sc_hd__a21oi_2 _19974_ (.A1(_09221_),
    .A2(_09217_),
    .B1(_09212_),
    .Y(_09680_));
 sky130_fd_sc_hd__o31ai_4 _19975_ (.A1(_08803_),
    .A2(_09216_),
    .A3(_09218_),
    .B1(_09213_),
    .Y(_09681_));
 sky130_fd_sc_hd__a21oi_1 _19976_ (.A1(_09213_),
    .A2(_09222_),
    .B1(_09679_),
    .Y(_09682_));
 sky130_fd_sc_hd__nand2_2 _19977_ (.A(_09678_),
    .B(_09681_),
    .Y(_09683_));
 sky130_fd_sc_hd__o221ai_4 _19978_ (.A1(net224),
    .A2(_09210_),
    .B1(_09672_),
    .B2(_09676_),
    .C1(_09222_),
    .Y(_09684_));
 sky130_fd_sc_hd__o22ai_2 _19979_ (.A1(_07691_),
    .A2(net371),
    .B1(_09681_),
    .B2(_09678_),
    .Y(_09685_));
 sky130_fd_sc_hd__nand3_1 _19980_ (.A(_09683_),
    .B(_09684_),
    .C(net354),
    .Y(_09687_));
 sky130_fd_sc_hd__o2bb2ai_4 _19981_ (.A1_N(_07724_),
    .A2_N(_09669_),
    .B1(_09682_),
    .B2(_09685_),
    .Y(_09688_));
 sky130_fd_sc_hd__a2bb2oi_2 _19982_ (.A1_N(_07242_),
    .A2_N(_07243_),
    .B1(_09671_),
    .B2(_09687_),
    .Y(_09689_));
 sky130_fd_sc_hd__o21ai_2 _19983_ (.A1(_07242_),
    .A2(_07243_),
    .B1(_09688_),
    .Y(_09690_));
 sky130_fd_sc_hd__o211a_1 _19984_ (.A1(_07244_),
    .A2(_07245_),
    .B1(_09671_),
    .C1(_09687_),
    .X(_09691_));
 sky130_fd_sc_hd__a311o_4 _19985_ (.A1(_09683_),
    .A2(_09684_),
    .A3(net354),
    .B1(net222),
    .C1(_09670_),
    .X(_09692_));
 sky130_fd_sc_hd__nand2_1 _19986_ (.A(_09231_),
    .B(_09237_),
    .Y(_09693_));
 sky130_fd_sc_hd__o22ai_1 _19987_ (.A1(net227),
    .A2(_09226_),
    .B1(_09239_),
    .B2(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__nand4_2 _19988_ (.A(_09229_),
    .B(_09244_),
    .C(_09690_),
    .D(_09692_),
    .Y(_09695_));
 sky130_fd_sc_hd__o21ai_1 _19989_ (.A1(_09689_),
    .A2(_09691_),
    .B1(_09694_),
    .Y(_09696_));
 sky130_fd_sc_hd__o211ai_4 _19990_ (.A1(_08678_),
    .A2(_08700_),
    .B1(_09695_),
    .C1(_09696_),
    .Y(_09698_));
 sky130_fd_sc_hd__a211o_1 _19991_ (.A1(_09671_),
    .A2(_09687_),
    .B1(_08678_),
    .C1(_08700_),
    .X(_09699_));
 sky130_fd_sc_hd__o211ai_2 _19992_ (.A1(_09689_),
    .A2(_09691_),
    .B1(_09229_),
    .C1(_09244_),
    .Y(_09700_));
 sky130_fd_sc_hd__nand3_1 _19993_ (.A(_09694_),
    .B(_09692_),
    .C(_09690_),
    .Y(_09701_));
 sky130_fd_sc_hd__o211ai_4 _19994_ (.A1(_08678_),
    .A2(_08700_),
    .B1(_09700_),
    .C1(_09701_),
    .Y(_09702_));
 sky130_fd_sc_hd__nand2_4 _19995_ (.A(_09699_),
    .B(_09702_),
    .Y(_09703_));
 sky130_fd_sc_hd__o21ai_2 _19996_ (.A1(net338),
    .A2(_09688_),
    .B1(_09698_),
    .Y(_09704_));
 sky130_fd_sc_hd__o211a_1 _19997_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_09699_),
    .C1(_09702_),
    .X(_09705_));
 sky130_fd_sc_hd__o211ai_2 _19998_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_09699_),
    .C1(_09702_),
    .Y(_09706_));
 sky130_fd_sc_hd__o211a_1 _19999_ (.A1(_09688_),
    .A2(net338),
    .B1(net225),
    .C1(_09698_),
    .X(_09707_));
 sky130_fd_sc_hd__o211ai_4 _20000_ (.A1(_09688_),
    .A2(net338),
    .B1(net225),
    .C1(_09698_),
    .Y(_09709_));
 sky130_fd_sc_hd__nand2_1 _20001_ (.A(_09706_),
    .B(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__and3_1 _20002_ (.A(_08048_),
    .B(_08432_),
    .C(_08433_),
    .X(_09711_));
 sky130_fd_sc_hd__nand4b_1 _20003_ (.A_N(_08057_),
    .B(_08845_),
    .C(_08847_),
    .D(_09711_),
    .Y(_09712_));
 sky130_fd_sc_hd__nand3_2 _20004_ (.A(_09255_),
    .B(_09711_),
    .C(_08848_),
    .Y(_09713_));
 sky130_fd_sc_hd__nor3_1 _20005_ (.A(_09712_),
    .B(_09256_),
    .C(_09254_),
    .Y(_09714_));
 sky130_fd_sc_hd__nand3b_4 _20006_ (.A_N(_09712_),
    .B(_09257_),
    .C(_09255_),
    .Y(_09715_));
 sky130_fd_sc_hd__o211a_1 _20007_ (.A1(_09261_),
    .A2(_09254_),
    .B1(_09257_),
    .C1(_09713_),
    .X(_09716_));
 sky130_fd_sc_hd__o211ai_4 _20008_ (.A1(_09261_),
    .A2(_09254_),
    .B1(_09257_),
    .C1(_09713_),
    .Y(_09717_));
 sky130_fd_sc_hd__a31o_2 _20009_ (.A1(_09257_),
    .A2(_09265_),
    .A3(_09713_),
    .B1(_09714_),
    .X(_09718_));
 sky130_fd_sc_hd__inv_2 _20010_ (.A(_09718_),
    .Y(_09720_));
 sky130_fd_sc_hd__a21oi_2 _20011_ (.A1(_09715_),
    .A2(_09717_),
    .B1(_09710_),
    .Y(_09721_));
 sky130_fd_sc_hd__a31o_1 _20012_ (.A1(_09710_),
    .A2(_09715_),
    .A3(_09717_),
    .B1(_09840_),
    .X(_09722_));
 sky130_fd_sc_hd__and3_1 _20013_ (.A(_09703_),
    .B(_09818_),
    .C(_09796_),
    .X(_09723_));
 sky130_fd_sc_hd__or3_2 _20014_ (.A(net351),
    .B(_09807_),
    .C(_09704_),
    .X(_09724_));
 sky130_fd_sc_hd__nand4_4 _20015_ (.A(_09706_),
    .B(_09709_),
    .C(_09715_),
    .D(_09717_),
    .Y(_09725_));
 sky130_fd_sc_hd__o22ai_4 _20016_ (.A1(_09705_),
    .A2(_09707_),
    .B1(_09714_),
    .B2(_09716_),
    .Y(_09726_));
 sky130_fd_sc_hd__nand3_2 _20017_ (.A(_09726_),
    .B(net336),
    .C(_09725_),
    .Y(_09727_));
 sky130_fd_sc_hd__o221a_2 _20018_ (.A1(net336),
    .A2(_09703_),
    .B1(_09721_),
    .B2(_09722_),
    .C1(_11079_),
    .X(_09728_));
 sky130_fd_sc_hd__a211o_2 _20019_ (.A1(_09724_),
    .A2(_09727_),
    .B1(_11046_),
    .C1(_11057_),
    .X(_09729_));
 sky130_fd_sc_hd__a311oi_4 _20020_ (.A1(_09726_),
    .A2(net336),
    .A3(_09725_),
    .B1(net232),
    .C1(_09723_),
    .Y(_09731_));
 sky130_fd_sc_hd__nand3_4 _20021_ (.A(_09727_),
    .B(net234),
    .C(_09724_),
    .Y(_09732_));
 sky130_fd_sc_hd__o221ai_4 _20022_ (.A1(net336),
    .A2(_09703_),
    .B1(_09721_),
    .B2(_09722_),
    .C1(net232),
    .Y(_09733_));
 sky130_fd_sc_hd__a21oi_1 _20023_ (.A1(net251),
    .A2(_09268_),
    .B1(_09278_),
    .Y(_09734_));
 sky130_fd_sc_hd__o22a_1 _20024_ (.A1(_09252_),
    .A2(_09273_),
    .B1(_09270_),
    .B2(_09278_),
    .X(_09735_));
 sky130_fd_sc_hd__o22ai_4 _20025_ (.A1(_09252_),
    .A2(_09273_),
    .B1(_09270_),
    .B2(_09278_),
    .Y(_09736_));
 sky130_fd_sc_hd__o2bb2ai_4 _20026_ (.A1_N(_09732_),
    .A2_N(_09733_),
    .B1(_09734_),
    .B2(_09274_),
    .Y(_09737_));
 sky130_fd_sc_hd__nand3_4 _20027_ (.A(_09735_),
    .B(_09733_),
    .C(_09732_),
    .Y(_09738_));
 sky130_fd_sc_hd__nand3_2 _20028_ (.A(_09737_),
    .B(_09738_),
    .C(net333),
    .Y(_09739_));
 sky130_fd_sc_hd__a21oi_1 _20029_ (.A1(_09293_),
    .A2(_09290_),
    .B1(_09287_),
    .Y(_09740_));
 sky130_fd_sc_hd__o21bai_2 _20030_ (.A1(_09289_),
    .A2(_09294_),
    .B1_N(_09287_),
    .Y(_09742_));
 sky130_fd_sc_hd__a31oi_4 _20031_ (.A1(_09737_),
    .A2(_09738_),
    .A3(net333),
    .B1(net251),
    .Y(_09743_));
 sky130_fd_sc_hd__a31o_1 _20032_ (.A1(_09737_),
    .A2(_09738_),
    .A3(net333),
    .B1(net251),
    .X(_09744_));
 sky130_fd_sc_hd__a311oi_4 _20033_ (.A1(_09737_),
    .A2(_09738_),
    .A3(net333),
    .B1(net251),
    .C1(_09728_),
    .Y(_09745_));
 sky130_fd_sc_hd__a311o_1 _20034_ (.A1(_09737_),
    .A2(_09738_),
    .A3(net333),
    .B1(net251),
    .C1(_09728_),
    .X(_09746_));
 sky130_fd_sc_hd__a2bb2oi_4 _20035_ (.A1_N(_06305_),
    .A2_N(net283),
    .B1(_09729_),
    .B2(_09739_),
    .Y(_09747_));
 sky130_fd_sc_hd__a22o_1 _20036_ (.A1(_06306_),
    .A2(_06308_),
    .B1(_09729_),
    .B2(_09739_),
    .X(_09748_));
 sky130_fd_sc_hd__nand3_2 _20037_ (.A(_09742_),
    .B(_09746_),
    .C(_09748_),
    .Y(_09749_));
 sky130_fd_sc_hd__o21ai_2 _20038_ (.A1(_09745_),
    .A2(_09747_),
    .B1(_09740_),
    .Y(_09750_));
 sky130_fd_sc_hd__a211o_2 _20039_ (.A1(_09729_),
    .A2(_09739_),
    .B1(_12670_),
    .C1(net327),
    .X(_09751_));
 sky130_fd_sc_hd__inv_2 _20040_ (.A(_09751_),
    .Y(_09753_));
 sky130_fd_sc_hd__o211a_1 _20041_ (.A1(_12670_),
    .A2(net327),
    .B1(_09749_),
    .C1(_09750_),
    .X(_09754_));
 sky130_fd_sc_hd__nand3_2 _20042_ (.A(_09749_),
    .B(_09750_),
    .C(net312),
    .Y(_09755_));
 sky130_fd_sc_hd__a31o_2 _20043_ (.A1(net312),
    .A2(_09749_),
    .A3(_09750_),
    .B1(_09753_),
    .X(_09756_));
 sky130_fd_sc_hd__a2bb2oi_1 _20044_ (.A1_N(_06009_),
    .A2_N(_06010_),
    .B1(_09751_),
    .B2(_09755_),
    .Y(_09757_));
 sky130_fd_sc_hd__o22ai_4 _20045_ (.A1(_06009_),
    .A2(_06010_),
    .B1(_09753_),
    .B2(_09754_),
    .Y(_09758_));
 sky130_fd_sc_hd__a31o_1 _20046_ (.A1(_09749_),
    .A2(_09750_),
    .A3(net312),
    .B1(net253),
    .X(_09759_));
 sky130_fd_sc_hd__o211a_1 _20047_ (.A1(net286),
    .A2(_06012_),
    .B1(_09751_),
    .C1(_09755_),
    .X(_09760_));
 sky130_fd_sc_hd__o211ai_4 _20048_ (.A1(net286),
    .A2(_06012_),
    .B1(_09751_),
    .C1(_09755_),
    .Y(_09761_));
 sky130_fd_sc_hd__nand2_1 _20049_ (.A(_09310_),
    .B(_09316_),
    .Y(_09762_));
 sky130_fd_sc_hd__nand3_1 _20050_ (.A(_09309_),
    .B(_09310_),
    .C(_09316_),
    .Y(_09764_));
 sky130_fd_sc_hd__o22ai_1 _20051_ (.A1(net262),
    .A2(_09301_),
    .B1(_09762_),
    .B2(_09308_),
    .Y(_09765_));
 sky130_fd_sc_hd__a31oi_4 _20052_ (.A1(_09309_),
    .A2(_09310_),
    .A3(_09316_),
    .B1(_09312_),
    .Y(_09766_));
 sky130_fd_sc_hd__o2111ai_4 _20053_ (.A1(_09308_),
    .A2(_09762_),
    .B1(_09761_),
    .C1(_09758_),
    .D1(_09314_),
    .Y(_09767_));
 sky130_fd_sc_hd__o21ai_1 _20054_ (.A1(_09757_),
    .A2(_09760_),
    .B1(_09765_),
    .Y(_09768_));
 sky130_fd_sc_hd__nand3_4 _20055_ (.A(_09767_),
    .B(_09768_),
    .C(net308),
    .Y(_09769_));
 sky130_fd_sc_hd__a211o_1 _20056_ (.A1(_09751_),
    .A2(_09755_),
    .B1(_00011_),
    .C1(net323),
    .X(_09770_));
 sky130_fd_sc_hd__o21ai_1 _20057_ (.A1(_09757_),
    .A2(_09760_),
    .B1(_09766_),
    .Y(_09771_));
 sky130_fd_sc_hd__o211ai_1 _20058_ (.A1(_09753_),
    .A2(_09759_),
    .B1(_09758_),
    .C1(_09765_),
    .Y(_09772_));
 sky130_fd_sc_hd__nand3_1 _20059_ (.A(_09772_),
    .B(net308),
    .C(_09771_),
    .Y(_09773_));
 sky130_fd_sc_hd__o21ai_2 _20060_ (.A1(net309),
    .A2(_09756_),
    .B1(_09769_),
    .Y(_09775_));
 sky130_fd_sc_hd__inv_2 _20061_ (.A(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__o311a_1 _20062_ (.A1(net308),
    .A2(_09753_),
    .A3(_09754_),
    .B1(_09769_),
    .C1(net261),
    .X(_09777_));
 sky130_fd_sc_hd__o211ai_4 _20063_ (.A1(net309),
    .A2(_09756_),
    .B1(_09769_),
    .C1(net261),
    .Y(_09778_));
 sky130_fd_sc_hd__o211ai_4 _20064_ (.A1(_05765_),
    .A2(net289),
    .B1(_09770_),
    .C1(_09773_),
    .Y(_09779_));
 sky130_fd_sc_hd__nand2_1 _20065_ (.A(_09778_),
    .B(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__and4_1 _20066_ (.A(_08124_),
    .B(_08126_),
    .C(_08509_),
    .D(_08511_),
    .X(_09781_));
 sky130_fd_sc_hd__nand3_2 _20067_ (.A(_09328_),
    .B(_09781_),
    .C(_08922_),
    .Y(_09782_));
 sky130_fd_sc_hd__o211ai_4 _20068_ (.A1(_09332_),
    .A2(_09327_),
    .B1(_09330_),
    .C1(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__inv_2 _20069_ (.A(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__and4_1 _20070_ (.A(_09781_),
    .B(_08921_),
    .C(_08919_),
    .D(_08128_),
    .X(_09786_));
 sky130_fd_sc_hd__nand3_4 _20071_ (.A(_09328_),
    .B(_09330_),
    .C(_09786_),
    .Y(_09787_));
 sky130_fd_sc_hd__inv_2 _20072_ (.A(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__a31o_1 _20073_ (.A1(_09330_),
    .A2(_09337_),
    .A3(_09782_),
    .B1(_09788_),
    .X(_09789_));
 sky130_fd_sc_hd__a21oi_2 _20074_ (.A1(_09783_),
    .A2(_09787_),
    .B1(_09780_),
    .Y(_09790_));
 sky130_fd_sc_hd__a31o_1 _20075_ (.A1(_09780_),
    .A2(_09783_),
    .A3(_09787_),
    .B1(_01973_),
    .X(_09791_));
 sky130_fd_sc_hd__o311a_2 _20076_ (.A1(net308),
    .A2(_09753_),
    .A3(_09754_),
    .B1(_09769_),
    .C1(_01973_),
    .X(_09792_));
 sky130_fd_sc_hd__or3_1 _20077_ (.A(_01940_),
    .B(net303),
    .C(_09775_),
    .X(_09793_));
 sky130_fd_sc_hd__nand4_4 _20078_ (.A(_09778_),
    .B(_09779_),
    .C(_09783_),
    .D(_09787_),
    .Y(_09794_));
 sky130_fd_sc_hd__a22o_1 _20079_ (.A1(_09778_),
    .A2(_09779_),
    .B1(_09783_),
    .B2(_09787_),
    .X(_09795_));
 sky130_fd_sc_hd__nand3_2 _20080_ (.A(_09795_),
    .B(net279),
    .C(_09794_),
    .Y(_09797_));
 sky130_fd_sc_hd__a31o_1 _20081_ (.A1(_09795_),
    .A2(net279),
    .A3(_09794_),
    .B1(_09792_),
    .X(_09798_));
 sky130_fd_sc_hd__o221a_2 _20082_ (.A1(net279),
    .A2(_09776_),
    .B1(_09790_),
    .B2(_09791_),
    .C1(_04040_),
    .X(_09799_));
 sky130_fd_sc_hd__a211o_2 _20083_ (.A1(_09793_),
    .A2(_09797_),
    .B1(_04008_),
    .C1(net300),
    .X(_09800_));
 sky130_fd_sc_hd__a311oi_4 _20084_ (.A1(_09795_),
    .A2(net279),
    .A3(_09794_),
    .B1(net291),
    .C1(_09792_),
    .Y(_09801_));
 sky130_fd_sc_hd__nand3_4 _20085_ (.A(_09797_),
    .B(net267),
    .C(_09793_),
    .Y(_09802_));
 sky130_fd_sc_hd__o221ai_4 _20086_ (.A1(net279),
    .A2(_09776_),
    .B1(_09790_),
    .B2(_09791_),
    .C1(net291),
    .Y(_09803_));
 sky130_fd_sc_hd__a21oi_1 _20087_ (.A1(net293),
    .A2(_09340_),
    .B1(_09343_),
    .Y(_09804_));
 sky130_fd_sc_hd__o32a_1 _20088_ (.A1(_05242_),
    .A2(net317),
    .A3(_09340_),
    .B1(_09343_),
    .B2(_09348_),
    .X(_09805_));
 sky130_fd_sc_hd__a21oi_1 _20089_ (.A1(_09347_),
    .A2(_09343_),
    .B1(_09348_),
    .Y(_09806_));
 sky130_fd_sc_hd__a21oi_1 _20090_ (.A1(_09802_),
    .A2(_09803_),
    .B1(_09805_),
    .Y(_09808_));
 sky130_fd_sc_hd__o2bb2ai_4 _20091_ (.A1_N(_09802_),
    .A2_N(_09803_),
    .B1(_09804_),
    .B2(_09345_),
    .Y(_09809_));
 sky130_fd_sc_hd__and3_1 _20092_ (.A(_09805_),
    .B(_09803_),
    .C(_09802_),
    .X(_09810_));
 sky130_fd_sc_hd__nand3_4 _20093_ (.A(_09805_),
    .B(_09803_),
    .C(_09802_),
    .Y(_09811_));
 sky130_fd_sc_hd__nand3_1 _20094_ (.A(_09809_),
    .B(_09811_),
    .C(net276),
    .Y(_09812_));
 sky130_fd_sc_hd__o22ai_1 _20095_ (.A1(_04008_),
    .A2(net300),
    .B1(_09808_),
    .B2(_09810_),
    .Y(_09813_));
 sky130_fd_sc_hd__a31oi_4 _20096_ (.A1(_09809_),
    .A2(_09811_),
    .A3(net276),
    .B1(_09799_),
    .Y(_09814_));
 sky130_fd_sc_hd__inv_2 _20097_ (.A(_09814_),
    .Y(_09815_));
 sky130_fd_sc_hd__o311a_1 _20098_ (.A1(_08553_),
    .A2(_08952_),
    .A3(_08954_),
    .B1(_09361_),
    .C1(_08950_),
    .X(_09816_));
 sky130_fd_sc_hd__and2_1 _20099_ (.A(_09362_),
    .B(_09365_),
    .X(_09817_));
 sky130_fd_sc_hd__nand2_1 _20100_ (.A(_09362_),
    .B(_09365_),
    .Y(_09819_));
 sky130_fd_sc_hd__o21ai_2 _20101_ (.A1(net299),
    .A2(_09359_),
    .B1(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__a31oi_2 _20102_ (.A1(_09809_),
    .A2(_09811_),
    .A3(net276),
    .B1(net293),
    .Y(_09821_));
 sky130_fd_sc_hd__a311oi_4 _20103_ (.A1(_09809_),
    .A2(_09811_),
    .A3(net276),
    .B1(net293),
    .C1(_09799_),
    .Y(_09822_));
 sky130_fd_sc_hd__a311o_1 _20104_ (.A1(_09809_),
    .A2(_09811_),
    .A3(net276),
    .B1(net293),
    .C1(_09799_),
    .X(_09823_));
 sky130_fd_sc_hd__a2bb2oi_4 _20105_ (.A1_N(_05242_),
    .A2_N(net317),
    .B1(_09800_),
    .B2(_09812_),
    .Y(_09824_));
 sky130_fd_sc_hd__o221ai_2 _20106_ (.A1(_05242_),
    .A2(net317),
    .B1(_09798_),
    .B2(net276),
    .C1(_09813_),
    .Y(_09825_));
 sky130_fd_sc_hd__o211ai_1 _20107_ (.A1(_09363_),
    .A2(_09816_),
    .B1(_09823_),
    .C1(_09825_),
    .Y(_09826_));
 sky130_fd_sc_hd__o22ai_1 _20108_ (.A1(_09360_),
    .A2(_09817_),
    .B1(_09822_),
    .B2(_09824_),
    .Y(_09827_));
 sky130_fd_sc_hd__nand3_1 _20109_ (.A(_09826_),
    .B(_09827_),
    .C(net273),
    .Y(_09828_));
 sky130_fd_sc_hd__or3_1 _20110_ (.A(net297),
    .B(_05232_),
    .C(_09814_),
    .X(_09830_));
 sky130_fd_sc_hd__o21ai_1 _20111_ (.A1(net295),
    .A2(_09814_),
    .B1(_09820_),
    .Y(_09831_));
 sky130_fd_sc_hd__o22ai_2 _20112_ (.A1(_09363_),
    .A2(_09816_),
    .B1(_09822_),
    .B2(_09824_),
    .Y(_09832_));
 sky130_fd_sc_hd__o221ai_4 _20113_ (.A1(net297),
    .A2(_05232_),
    .B1(_09822_),
    .B2(_09831_),
    .C1(_09832_),
    .Y(_09833_));
 sky130_fd_sc_hd__o21ai_2 _20114_ (.A1(net273),
    .A2(_09814_),
    .B1(_09833_),
    .Y(_09834_));
 sky130_fd_sc_hd__o211a_1 _20115_ (.A1(_09815_),
    .A2(net273),
    .B1(net298),
    .C1(_09828_),
    .X(_09835_));
 sky130_fd_sc_hd__o211ai_2 _20116_ (.A1(_09815_),
    .A2(net273),
    .B1(net298),
    .C1(_09828_),
    .Y(_09836_));
 sky130_fd_sc_hd__and3_1 _20117_ (.A(_09833_),
    .B(net299),
    .C(_09830_),
    .X(_09837_));
 sky130_fd_sc_hd__o211ai_4 _20118_ (.A1(net273),
    .A2(_09814_),
    .B1(net299),
    .C1(_09833_),
    .Y(_09838_));
 sky130_fd_sc_hd__a21oi_1 _20119_ (.A1(_09383_),
    .A2(_09384_),
    .B1(_09374_),
    .Y(_09839_));
 sky130_fd_sc_hd__a22o_1 _20120_ (.A1(_02148_),
    .A2(_09373_),
    .B1(_09383_),
    .B2(_09384_),
    .X(_09841_));
 sky130_fd_sc_hd__o2bb2ai_1 _20121_ (.A1_N(_09836_),
    .A2_N(_09838_),
    .B1(_09839_),
    .B2(_09376_),
    .Y(_09842_));
 sky130_fd_sc_hd__nand4_1 _20122_ (.A(_09377_),
    .B(_09836_),
    .C(_09838_),
    .D(_09841_),
    .Y(_09843_));
 sky130_fd_sc_hd__a22o_1 _20123_ (.A1(_05482_),
    .A2(_05484_),
    .B1(_09842_),
    .B2(_09843_),
    .X(_09844_));
 sky130_fd_sc_hd__a211o_2 _20124_ (.A1(_09830_),
    .A2(_09833_),
    .B1(_05481_),
    .C1(_05483_),
    .X(_09845_));
 sky130_fd_sc_hd__nand3_2 _20125_ (.A(_09842_),
    .B(_09843_),
    .C(net246),
    .Y(_09846_));
 sky130_fd_sc_hd__nand2_1 _20126_ (.A(_09845_),
    .B(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__or3_1 _20127_ (.A(net266),
    .B(_05751_),
    .C(_09847_),
    .X(_09848_));
 sky130_fd_sc_hd__a2bb2oi_1 _20128_ (.A1_N(_02049_),
    .A2_N(net343),
    .B1(_09845_),
    .B2(_09846_),
    .Y(_09849_));
 sky130_fd_sc_hd__o221ai_4 _20129_ (.A1(_02049_),
    .A2(_02071_),
    .B1(net246),
    .B2(_09834_),
    .C1(_09844_),
    .Y(_09850_));
 sky130_fd_sc_hd__o211a_2 _20130_ (.A1(_02093_),
    .A2(_02115_),
    .B1(_09845_),
    .C1(_09846_),
    .X(_09852_));
 sky130_fd_sc_hd__o211ai_2 _20131_ (.A1(_02093_),
    .A2(_02115_),
    .B1(_09845_),
    .C1(_09846_),
    .Y(_09853_));
 sky130_fd_sc_hd__o22a_1 _20132_ (.A1(_09395_),
    .A2(_09389_),
    .B1(_09399_),
    .B2(_09397_),
    .X(_09854_));
 sky130_fd_sc_hd__o22ai_4 _20133_ (.A1(_09395_),
    .A2(_09389_),
    .B1(_09399_),
    .B2(_09397_),
    .Y(_09855_));
 sky130_fd_sc_hd__a31o_1 _20134_ (.A1(_02137_),
    .A2(_09845_),
    .A3(_09846_),
    .B1(_09855_),
    .X(_09856_));
 sky130_fd_sc_hd__nand3_2 _20135_ (.A(_09850_),
    .B(_09854_),
    .C(_09853_),
    .Y(_09857_));
 sky130_fd_sc_hd__o21ai_2 _20136_ (.A1(_09849_),
    .A2(_09852_),
    .B1(_09855_),
    .Y(_09858_));
 sky130_fd_sc_hd__nand3_1 _20137_ (.A(_09850_),
    .B(_09853_),
    .C(_09855_),
    .Y(_09859_));
 sky130_fd_sc_hd__o21ai_1 _20138_ (.A1(_09849_),
    .A2(_09852_),
    .B1(_09854_),
    .Y(_09860_));
 sky130_fd_sc_hd__nand3_2 _20139_ (.A(_09860_),
    .B(net242),
    .C(_09859_),
    .Y(_09861_));
 sky130_fd_sc_hd__o311a_1 _20140_ (.A1(_05481_),
    .A2(_05483_),
    .A3(_09834_),
    .B1(_09844_),
    .C1(_05754_),
    .X(_09863_));
 sky130_fd_sc_hd__a211o_1 _20141_ (.A1(_09845_),
    .A2(_09846_),
    .B1(net266),
    .C1(_05751_),
    .X(_09864_));
 sky130_fd_sc_hd__nand3_1 _20142_ (.A(_09858_),
    .B(net242),
    .C(_09857_),
    .Y(_09865_));
 sky130_fd_sc_hd__o21ai_2 _20143_ (.A1(net241),
    .A2(_09847_),
    .B1(_09861_),
    .Y(_09866_));
 sky130_fd_sc_hd__inv_2 _20144_ (.A(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__and3_1 _20145_ (.A(_09861_),
    .B(_05995_),
    .C(_09848_),
    .X(_09868_));
 sky130_fd_sc_hd__or3_1 _20146_ (.A(net259),
    .B(net257),
    .C(_09866_),
    .X(_09869_));
 sky130_fd_sc_hd__a311oi_4 _20147_ (.A1(_09858_),
    .A2(net242),
    .A3(_09857_),
    .B1(_09863_),
    .C1(_00251_),
    .Y(_09870_));
 sky130_fd_sc_hd__nand3_4 _20148_ (.A(_09865_),
    .B(net320),
    .C(_09864_),
    .Y(_09871_));
 sky130_fd_sc_hd__o311a_1 _20149_ (.A1(net266),
    .A2(_05751_),
    .A3(_09847_),
    .B1(_09861_),
    .C1(_00251_),
    .X(_09872_));
 sky130_fd_sc_hd__o211ai_4 _20150_ (.A1(_00174_),
    .A2(net344),
    .B1(_09848_),
    .C1(_09861_),
    .Y(_09874_));
 sky130_fd_sc_hd__a21oi_1 _20151_ (.A1(net326),
    .A2(_09408_),
    .B1(_09413_),
    .Y(_09875_));
 sky130_fd_sc_hd__a21oi_2 _20152_ (.A1(_09415_),
    .A2(_09394_),
    .B1(_09414_),
    .Y(_09876_));
 sky130_fd_sc_hd__o21ai_1 _20153_ (.A1(_09414_),
    .A2(_09416_),
    .B1(_09419_),
    .Y(_09877_));
 sky130_fd_sc_hd__a21oi_2 _20154_ (.A1(_09417_),
    .A2(_09413_),
    .B1(_09418_),
    .Y(_09878_));
 sky130_fd_sc_hd__a21oi_1 _20155_ (.A1(_09871_),
    .A2(_09874_),
    .B1(_09877_),
    .Y(_09879_));
 sky130_fd_sc_hd__o2bb2ai_4 _20156_ (.A1_N(_09871_),
    .A2_N(_09874_),
    .B1(_09875_),
    .B2(_09416_),
    .Y(_09880_));
 sky130_fd_sc_hd__o211a_1 _20157_ (.A1(_09418_),
    .A2(_09876_),
    .B1(_09874_),
    .C1(_09871_),
    .X(_09881_));
 sky130_fd_sc_hd__o211ai_4 _20158_ (.A1(_09418_),
    .A2(_09876_),
    .B1(_09874_),
    .C1(_09871_),
    .Y(_09882_));
 sky130_fd_sc_hd__a31oi_2 _20159_ (.A1(_09877_),
    .A2(_09874_),
    .A3(_09871_),
    .B1(_05995_),
    .Y(_09883_));
 sky130_fd_sc_hd__o211ai_4 _20160_ (.A1(net259),
    .A2(net257),
    .B1(_09880_),
    .C1(_09882_),
    .Y(_09884_));
 sky130_fd_sc_hd__o22ai_2 _20161_ (.A1(net259),
    .A2(net257),
    .B1(_09879_),
    .B2(_09881_),
    .Y(_09885_));
 sky130_fd_sc_hd__a31o_1 _20162_ (.A1(net240),
    .A2(_09880_),
    .A3(_09882_),
    .B1(_09868_),
    .X(_09886_));
 sky130_fd_sc_hd__a31oi_4 _20163_ (.A1(_11309_),
    .A2(_09409_),
    .A3(_09422_),
    .B1(_09436_),
    .Y(_09887_));
 sky130_fd_sc_hd__a31oi_4 _20164_ (.A1(_11298_),
    .A2(_09424_),
    .A3(_09427_),
    .B1(_09437_),
    .Y(_09888_));
 sky130_fd_sc_hd__a211oi_4 _20165_ (.A1(_09883_),
    .A2(_09880_),
    .B1(_09868_),
    .C1(net326),
    .Y(_09889_));
 sky130_fd_sc_hd__o221ai_4 _20166_ (.A1(_12867_),
    .A2(_12877_),
    .B1(net240),
    .B2(_09866_),
    .C1(_09884_),
    .Y(_09890_));
 sky130_fd_sc_hd__a2bb2oi_2 _20167_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_09869_),
    .B2(_09884_),
    .Y(_09891_));
 sky130_fd_sc_hd__o211ai_4 _20168_ (.A1(_09867_),
    .A2(net240),
    .B1(net326),
    .C1(_09885_),
    .Y(_09892_));
 sky130_fd_sc_hd__o211ai_1 _20169_ (.A1(_09432_),
    .A2(_09887_),
    .B1(_09890_),
    .C1(_09892_),
    .Y(_09893_));
 sky130_fd_sc_hd__o22ai_1 _20170_ (.A1(_09430_),
    .A2(_09888_),
    .B1(_09889_),
    .B2(_09891_),
    .Y(_09895_));
 sky130_fd_sc_hd__nand3_2 _20171_ (.A(_09895_),
    .B(net212),
    .C(_09893_),
    .Y(_09896_));
 sky130_fd_sc_hd__o221a_1 _20172_ (.A1(_06286_),
    .A2(_06288_),
    .B1(_09867_),
    .B2(net240),
    .C1(_09885_),
    .X(_09897_));
 sky130_fd_sc_hd__a22o_1 _20173_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_09869_),
    .B2(_09884_),
    .X(_09898_));
 sky130_fd_sc_hd__o211ai_4 _20174_ (.A1(_09430_),
    .A2(_09888_),
    .B1(_09890_),
    .C1(_09892_),
    .Y(_09899_));
 sky130_fd_sc_hd__o22ai_4 _20175_ (.A1(_09432_),
    .A2(_09887_),
    .B1(_09889_),
    .B2(_09891_),
    .Y(_09900_));
 sky130_fd_sc_hd__o211ai_2 _20176_ (.A1(_06291_),
    .A2(_06292_),
    .B1(_09899_),
    .C1(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__a31oi_4 _20177_ (.A1(_09900_),
    .A2(net212),
    .A3(_09899_),
    .B1(_09897_),
    .Y(_09902_));
 sky130_fd_sc_hd__o211a_1 _20178_ (.A1(_09886_),
    .A2(net212),
    .B1(_11309_),
    .C1(_09896_),
    .X(_09903_));
 sky130_fd_sc_hd__o211ai_4 _20179_ (.A1(_09886_),
    .A2(net212),
    .B1(_11309_),
    .C1(_09896_),
    .Y(_09904_));
 sky130_fd_sc_hd__o211ai_4 _20180_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_09898_),
    .C1(_09901_),
    .Y(_09906_));
 sky130_fd_sc_hd__inv_2 _20181_ (.A(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__a21oi_1 _20182_ (.A1(_09446_),
    .A2(_10025_),
    .B1(_09454_),
    .Y(_09908_));
 sky130_fd_sc_hd__a21o_1 _20183_ (.A1(_09451_),
    .A2(_09454_),
    .B1(_09448_),
    .X(_09909_));
 sky130_fd_sc_hd__a21oi_1 _20184_ (.A1(_09904_),
    .A2(_09906_),
    .B1(_09909_),
    .Y(_09910_));
 sky130_fd_sc_hd__o2bb2ai_1 _20185_ (.A1_N(_09904_),
    .A2_N(_09906_),
    .B1(_09908_),
    .B2(_09450_),
    .Y(_09911_));
 sky130_fd_sc_hd__o211ai_2 _20186_ (.A1(_09448_),
    .A2(_09457_),
    .B1(_09904_),
    .C1(_09906_),
    .Y(_09912_));
 sky130_fd_sc_hd__o21ai_1 _20187_ (.A1(_06608_),
    .A2(net237),
    .B1(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__nand3_4 _20188_ (.A(_09911_),
    .B(_09912_),
    .C(net211),
    .Y(_09914_));
 sky130_fd_sc_hd__or3_1 _20189_ (.A(_06608_),
    .B(net237),
    .C(_09902_),
    .X(_09915_));
 sky130_fd_sc_hd__o32a_1 _20190_ (.A1(_06608_),
    .A2(net237),
    .A3(_09902_),
    .B1(_09910_),
    .B2(_09913_),
    .X(_09917_));
 sky130_fd_sc_hd__o21ai_2 _20191_ (.A1(net211),
    .A2(_09902_),
    .B1(_09914_),
    .Y(_09918_));
 sky130_fd_sc_hd__a21oi_2 _20192_ (.A1(_09914_),
    .A2(_09915_),
    .B1(_10015_),
    .Y(_09919_));
 sky130_fd_sc_hd__a22o_1 _20193_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_09914_),
    .B2(_09915_),
    .X(_09920_));
 sky130_fd_sc_hd__o221a_1 _20194_ (.A1(net365),
    .A2(net364),
    .B1(net211),
    .B2(_09902_),
    .C1(_09914_),
    .X(_09921_));
 sky130_fd_sc_hd__o221ai_4 _20195_ (.A1(net365),
    .A2(net364),
    .B1(net211),
    .B2(_09902_),
    .C1(_09914_),
    .Y(_09922_));
 sky130_fd_sc_hd__a21oi_1 _20196_ (.A1(_09920_),
    .A2(_09922_),
    .B1(_09585_),
    .Y(_09923_));
 sky130_fd_sc_hd__o21ai_2 _20197_ (.A1(_09919_),
    .A2(_09921_),
    .B1(_09584_),
    .Y(_09924_));
 sky130_fd_sc_hd__o21ai_1 _20198_ (.A1(_09465_),
    .A2(_09583_),
    .B1(_09922_),
    .Y(_09925_));
 sky130_fd_sc_hd__o221ai_4 _20199_ (.A1(_09465_),
    .A2(_09583_),
    .B1(_09918_),
    .B2(_10025_),
    .C1(_09920_),
    .Y(_09926_));
 sky130_fd_sc_hd__o22ai_1 _20200_ (.A1(net230),
    .A2(_06901_),
    .B1(_09919_),
    .B2(_09925_),
    .Y(_09928_));
 sky130_fd_sc_hd__nand3_1 _20201_ (.A(_09924_),
    .B(_09926_),
    .C(net208),
    .Y(_09929_));
 sky130_fd_sc_hd__and3_1 _20202_ (.A(_06900_),
    .B(_06902_),
    .C(_09918_),
    .X(_09930_));
 sky130_fd_sc_hd__or3_1 _20203_ (.A(net230),
    .B(_06901_),
    .C(_09917_),
    .X(_09931_));
 sky130_fd_sc_hd__o21ai_2 _20204_ (.A1(_09923_),
    .A2(_09928_),
    .B1(_09931_),
    .Y(_09932_));
 sky130_fd_sc_hd__inv_2 _20205_ (.A(_09932_),
    .Y(_09933_));
 sky130_fd_sc_hd__o21a_1 _20206_ (.A1(_07888_),
    .A2(_09473_),
    .B1(_09477_),
    .X(_09934_));
 sky130_fd_sc_hd__o21ai_1 _20207_ (.A1(_09477_),
    .A2(_09479_),
    .B1(_09482_),
    .Y(_09935_));
 sky130_fd_sc_hd__a311oi_2 _20208_ (.A1(_09924_),
    .A2(_09926_),
    .A3(net208),
    .B1(_09930_),
    .C1(_08918_),
    .Y(_09936_));
 sky130_fd_sc_hd__a311o_1 _20209_ (.A1(_09924_),
    .A2(_09926_),
    .A3(net208),
    .B1(_09930_),
    .C1(_08918_),
    .X(_09937_));
 sky130_fd_sc_hd__a21oi_1 _20210_ (.A1(_09929_),
    .A2(_09931_),
    .B1(_08907_),
    .Y(_09939_));
 sky130_fd_sc_hd__o21ai_1 _20211_ (.A1(_08819_),
    .A2(_08841_),
    .B1(_09932_),
    .Y(_09940_));
 sky130_fd_sc_hd__o211a_1 _20212_ (.A1(_09479_),
    .A2(_09934_),
    .B1(_09937_),
    .C1(_09940_),
    .X(_09941_));
 sky130_fd_sc_hd__o21ai_1 _20213_ (.A1(_09936_),
    .A2(_09939_),
    .B1(_09935_),
    .Y(_09942_));
 sky130_fd_sc_hd__o21ai_1 _20214_ (.A1(_07227_),
    .A2(net203),
    .B1(_09942_),
    .Y(_09943_));
 sky130_fd_sc_hd__a211o_1 _20215_ (.A1(_09929_),
    .A2(_09931_),
    .B1(_07227_),
    .C1(net203),
    .X(_09944_));
 sky130_fd_sc_hd__nand3_1 _20216_ (.A(_09940_),
    .B(_09935_),
    .C(_09937_),
    .Y(_09945_));
 sky130_fd_sc_hd__o22ai_2 _20217_ (.A1(_09479_),
    .A2(_09934_),
    .B1(_09936_),
    .B2(_09939_),
    .Y(_09946_));
 sky130_fd_sc_hd__o211ai_4 _20218_ (.A1(_07227_),
    .A2(net203),
    .B1(_09945_),
    .C1(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__o22a_1 _20219_ (.A1(net185),
    .A2(_09932_),
    .B1(_09941_),
    .B2(_09943_),
    .X(_09948_));
 sky130_fd_sc_hd__inv_2 _20220_ (.A(_09948_),
    .Y(_09950_));
 sky130_fd_sc_hd__o221a_1 _20221_ (.A1(net368),
    .A2(_07866_),
    .B1(net185),
    .B2(_09933_),
    .C1(_09947_),
    .X(_09951_));
 sky130_fd_sc_hd__o221ai_4 _20222_ (.A1(net368),
    .A2(_07866_),
    .B1(net185),
    .B2(_09933_),
    .C1(_09947_),
    .Y(_09952_));
 sky130_fd_sc_hd__a21oi_2 _20223_ (.A1(_09944_),
    .A2(_09947_),
    .B1(_07888_),
    .Y(_09953_));
 sky130_fd_sc_hd__o221ai_1 _20224_ (.A1(net185),
    .A2(_09932_),
    .B1(_09941_),
    .B2(_09943_),
    .C1(_07899_),
    .Y(_09954_));
 sky130_fd_sc_hd__a21oi_1 _20225_ (.A1(_09497_),
    .A2(_09581_),
    .B1(_09951_),
    .Y(_09955_));
 sky130_fd_sc_hd__nand3_1 _20226_ (.A(_09582_),
    .B(_09952_),
    .C(_09954_),
    .Y(_09956_));
 sky130_fd_sc_hd__o22ai_2 _20227_ (.A1(_09494_),
    .A2(_09580_),
    .B1(_09951_),
    .B2(_09953_),
    .Y(_09957_));
 sky130_fd_sc_hd__and3_1 _20228_ (.A(_09948_),
    .B(_07547_),
    .C(_07545_),
    .X(_09958_));
 sky130_fd_sc_hd__a211o_2 _20229_ (.A1(_09944_),
    .A2(_09947_),
    .B1(_07544_),
    .C1(net184),
    .X(_09959_));
 sky130_fd_sc_hd__nand3_2 _20230_ (.A(_09957_),
    .B(net163),
    .C(_09956_),
    .Y(_09961_));
 sky130_fd_sc_hd__a21oi_4 _20231_ (.A1(_09959_),
    .A2(_09961_),
    .B1(net160),
    .Y(_09962_));
 sky130_fd_sc_hd__inv_2 _20232_ (.A(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__o32a_1 _20233_ (.A1(net381),
    .A2(_06310_),
    .A3(_09505_),
    .B1(_09509_),
    .B2(_09512_),
    .X(_09964_));
 sky130_fd_sc_hd__a31o_1 _20234_ (.A1(_09957_),
    .A2(net163),
    .A3(_09956_),
    .B1(_07044_),
    .X(_09965_));
 sky130_fd_sc_hd__o221a_2 _20235_ (.A1(_06989_),
    .A2(net375),
    .B1(net163),
    .B2(_09950_),
    .C1(_09961_),
    .X(_09966_));
 sky130_fd_sc_hd__a21oi_2 _20236_ (.A1(_09959_),
    .A2(_09961_),
    .B1(_07033_),
    .Y(_09967_));
 sky130_fd_sc_hd__a22o_2 _20237_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_09959_),
    .B2(_09961_),
    .X(_09968_));
 sky130_fd_sc_hd__o221ai_4 _20238_ (.A1(_09507_),
    .A2(_09516_),
    .B1(_09958_),
    .B2(_09965_),
    .C1(_09968_),
    .Y(_09969_));
 sky130_fd_sc_hd__o21ai_2 _20239_ (.A1(_09966_),
    .A2(_09967_),
    .B1(_09964_),
    .Y(_09970_));
 sky130_fd_sc_hd__nand3_1 _20240_ (.A(_09970_),
    .B(net160),
    .C(_09969_),
    .Y(_09972_));
 sky130_fd_sc_hd__a31oi_4 _20241_ (.A1(_09970_),
    .A2(net160),
    .A3(_09969_),
    .B1(_09962_),
    .Y(_09973_));
 sky130_fd_sc_hd__a2bb2oi_1 _20242_ (.A1_N(net394),
    .A2_N(_06267_),
    .B1(_09963_),
    .B2(_09972_),
    .Y(_09974_));
 sky130_fd_sc_hd__a22o_1 _20243_ (.A1(_06256_),
    .A2(_06278_),
    .B1(_09963_),
    .B2(_09972_),
    .X(_09975_));
 sky130_fd_sc_hd__a31o_1 _20244_ (.A1(_09970_),
    .A2(net160),
    .A3(_09969_),
    .B1(_06343_),
    .X(_09976_));
 sky130_fd_sc_hd__o211a_1 _20245_ (.A1(net381),
    .A2(_06310_),
    .B1(_09963_),
    .C1(_09972_),
    .X(_09977_));
 sky130_fd_sc_hd__a31o_1 _20246_ (.A1(_09506_),
    .A2(_09518_),
    .A3(_09525_),
    .B1(_09523_),
    .X(_09978_));
 sky130_fd_sc_hd__a31oi_2 _20247_ (.A1(_09506_),
    .A2(_09518_),
    .A3(_09525_),
    .B1(_09523_),
    .Y(_09979_));
 sky130_fd_sc_hd__o21ai_2 _20248_ (.A1(_09974_),
    .A2(_09977_),
    .B1(_09978_),
    .Y(_09980_));
 sky130_fd_sc_hd__a21oi_1 _20249_ (.A1(_06332_),
    .A2(_09973_),
    .B1(_09978_),
    .Y(_09981_));
 sky130_fd_sc_hd__o211ai_4 _20250_ (.A1(_09962_),
    .A2(_09976_),
    .B1(_09979_),
    .C1(_09975_),
    .Y(_09983_));
 sky130_fd_sc_hd__nand3_2 _20251_ (.A(_09980_),
    .B(_09983_),
    .C(_08300_),
    .Y(_09984_));
 sky130_fd_sc_hd__a22oi_4 _20252_ (.A1(_08297_),
    .A2(_08299_),
    .B1(_09980_),
    .B2(_09983_),
    .Y(_09985_));
 sky130_fd_sc_hd__a311o_1 _20253_ (.A1(_09970_),
    .A2(net160),
    .A3(_09969_),
    .B1(_08300_),
    .C1(_09962_),
    .X(_09986_));
 sky130_fd_sc_hd__inv_2 _20254_ (.A(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__o21ai_2 _20255_ (.A1(_08300_),
    .A2(_09973_),
    .B1(_09984_),
    .Y(_09988_));
 sky130_fd_sc_hd__o211ai_4 _20256_ (.A1(_05556_),
    .A2(_09531_),
    .B1(_09530_),
    .C1(_09528_),
    .Y(_09989_));
 sky130_fd_sc_hd__nand2_1 _20257_ (.A(_09532_),
    .B(_09989_),
    .Y(_09990_));
 sky130_fd_sc_hd__o211ai_4 _20258_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_09532_),
    .C1(_09989_),
    .Y(_09991_));
 sky130_fd_sc_hd__a22o_1 _20259_ (.A1(net395),
    .A2(_05796_),
    .B1(_09532_),
    .B2(_09989_),
    .X(_09992_));
 sky130_fd_sc_hd__o211ai_4 _20260_ (.A1(net158),
    .A2(_08712_),
    .B1(_09991_),
    .C1(_09992_),
    .Y(_09994_));
 sky130_fd_sc_hd__o211ai_4 _20261_ (.A1(_08300_),
    .A2(_09973_),
    .B1(_09984_),
    .C1(_09994_),
    .Y(_09995_));
 sky130_fd_sc_hd__o311a_1 _20262_ (.A1(net180),
    .A2(_08298_),
    .A3(_09973_),
    .B1(_05851_),
    .C1(_09984_),
    .X(_09996_));
 sky130_fd_sc_hd__o31a_1 _20263_ (.A1(_09994_),
    .A2(_09987_),
    .A3(_09985_),
    .B1(_09995_),
    .X(_09997_));
 sky130_fd_sc_hd__o31ai_1 _20264_ (.A1(_09994_),
    .A2(_09987_),
    .A3(_09985_),
    .B1(_09995_),
    .Y(_09998_));
 sky130_fd_sc_hd__o22ai_4 _20265_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_09540_),
    .B2(_09543_),
    .Y(_09999_));
 sky130_fd_sc_hd__o2111ai_4 _20266_ (.A1(_03399_),
    .A2(_05491_),
    .B1(net396),
    .C1(_09541_),
    .D1(_09545_),
    .Y(_10000_));
 sky130_fd_sc_hd__o211ai_1 _20267_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_09999_),
    .C1(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__nand4_4 _20268_ (.A(_09997_),
    .B(_09999_),
    .C(_10000_),
    .D(_09125_),
    .Y(_10002_));
 sky130_fd_sc_hd__nand2_2 _20269_ (.A(_09998_),
    .B(_10001_),
    .Y(_10003_));
 sky130_fd_sc_hd__a21o_1 _20270_ (.A1(_10002_),
    .A2(_10003_),
    .B1(net143),
    .X(_10005_));
 sky130_fd_sc_hd__a21oi_2 _20271_ (.A1(_10002_),
    .A2(_10003_),
    .B1(_05239_),
    .Y(_10006_));
 sky130_fd_sc_hd__a21o_1 _20272_ (.A1(_10002_),
    .A2(_10003_),
    .B1(_05239_),
    .X(_10007_));
 sky130_fd_sc_hd__nand4_2 _20273_ (.A(_05207_),
    .B(_05229_),
    .C(_10002_),
    .D(_10003_),
    .Y(_10008_));
 sky130_fd_sc_hd__a31oi_1 _20274_ (.A1(_05239_),
    .A2(_10002_),
    .A3(_10003_),
    .B1(_09549_),
    .Y(_10009_));
 sky130_fd_sc_hd__a22oi_1 _20275_ (.A1(net1),
    .A2(_09548_),
    .B1(_10007_),
    .B2(_10008_),
    .Y(_10010_));
 sky130_fd_sc_hd__a21oi_1 _20276_ (.A1(_10007_),
    .A2(_10009_),
    .B1(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__o21a_1 _20277_ (.A1(_09562_),
    .A2(_10011_),
    .B1(_10005_),
    .X(_10012_));
 sky130_fd_sc_hd__nand2_1 _20278_ (.A(net1),
    .B(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__xor2_1 _20279_ (.A(net1),
    .B(_10012_),
    .X(_10014_));
 sky130_fd_sc_hd__and3_1 _20280_ (.A(_10014_),
    .B(_09577_),
    .C(_09575_),
    .X(_10016_));
 sky130_fd_sc_hd__a21oi_2 _20281_ (.A1(_09578_),
    .A2(_10012_),
    .B1(_10016_),
    .Y(_10017_));
 sky130_fd_sc_hd__xnor2_1 _20282_ (.A(_09569_),
    .B(_10017_),
    .Y(net84));
 sky130_fd_sc_hd__a31o_1 _20283_ (.A1(_09130_),
    .A2(_09565_),
    .A3(_10017_),
    .B1(_05051_),
    .X(_10018_));
 sky130_fd_sc_hd__o21ai_2 _20284_ (.A1(_09977_),
    .A2(_09978_),
    .B1(_09975_),
    .Y(_10019_));
 sky130_fd_sc_hd__or4_4 _20285_ (.A(net18),
    .B(net19),
    .C(net20),
    .D(_08723_),
    .X(_10020_));
 sky130_fd_sc_hd__and3b_4 _20286_ (.A_N(net21),
    .B(_10020_),
    .C(net410),
    .X(_10021_));
 sky130_fd_sc_hd__a21boi_4 _20287_ (.A1(_10020_),
    .A2(net410),
    .B1_N(net21),
    .Y(_10022_));
 sky130_fd_sc_hd__a21oi_4 _20288_ (.A1(_10020_),
    .A2(net410),
    .B1(net21),
    .Y(_10023_));
 sky130_fd_sc_hd__o311a_4 _20289_ (.A1(net19),
    .A2(net20),
    .A3(_09133_),
    .B1(net21),
    .C1(net410),
    .X(_10024_));
 sky130_fd_sc_hd__nor2_8 _20290_ (.A(_10021_),
    .B(_10022_),
    .Y(_10026_));
 sky130_fd_sc_hd__nor2_8 _20291_ (.A(net167),
    .B(_10024_),
    .Y(_10027_));
 sky130_fd_sc_hd__o21a_1 _20292_ (.A1(net170),
    .A2(net169),
    .B1(net33),
    .X(_10028_));
 sky130_fd_sc_hd__or3_1 _20293_ (.A(_10024_),
    .B(_03178_),
    .C(_10023_),
    .X(_10029_));
 sky130_fd_sc_hd__o221a_1 _20294_ (.A1(_05130_),
    .A2(_05152_),
    .B1(net170),
    .B2(net169),
    .C1(net33),
    .X(_10030_));
 sky130_fd_sc_hd__or3_1 _20295_ (.A(_09588_),
    .B(_09590_),
    .C(_10028_),
    .X(_10031_));
 sky130_fd_sc_hd__o41ai_4 _20296_ (.A1(_03178_),
    .A2(_09592_),
    .A3(_09593_),
    .A4(net153),
    .B1(_10031_),
    .Y(_10032_));
 sky130_fd_sc_hd__inv_2 _20297_ (.A(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__a22oi_2 _20298_ (.A1(_09141_),
    .A2(_09595_),
    .B1(_09601_),
    .B2(_09600_),
    .Y(_10034_));
 sky130_fd_sc_hd__a22o_1 _20299_ (.A1(_09141_),
    .A2(_09595_),
    .B1(_09601_),
    .B2(_09600_),
    .X(_10035_));
 sky130_fd_sc_hd__nand2_1 _20300_ (.A(_10035_),
    .B(_10033_),
    .Y(_10037_));
 sky130_fd_sc_hd__a221o_1 _20301_ (.A1(_09141_),
    .A2(_09595_),
    .B1(_09601_),
    .B2(_09600_),
    .C1(_10033_),
    .X(_10038_));
 sky130_fd_sc_hd__a21o_1 _20302_ (.A1(_10037_),
    .A2(_10038_),
    .B1(_05185_),
    .X(_10039_));
 sky130_fd_sc_hd__o21ai_2 _20303_ (.A1(net405),
    .A2(_10028_),
    .B1(_10039_),
    .Y(_10040_));
 sky130_fd_sc_hd__inv_2 _20304_ (.A(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__or3_2 _20305_ (.A(_05348_),
    .B(net401),
    .C(_10040_),
    .X(_10042_));
 sky130_fd_sc_hd__a311o_2 _20306_ (.A1(_10037_),
    .A2(_10038_),
    .A3(net405),
    .B1(net173),
    .C1(_10030_),
    .X(_10043_));
 sky130_fd_sc_hd__o221ai_4 _20307_ (.A1(_09134_),
    .A2(_09135_),
    .B1(_10028_),
    .B2(net405),
    .C1(_10039_),
    .Y(_10044_));
 sky130_fd_sc_hd__and2_1 _20308_ (.A(_10043_),
    .B(_10044_),
    .X(_10045_));
 sky130_fd_sc_hd__nand2_1 _20309_ (.A(_10043_),
    .B(_10044_),
    .Y(_10046_));
 sky130_fd_sc_hd__o21ai_2 _20310_ (.A1(_09612_),
    .A2(_09616_),
    .B1(_09610_),
    .Y(_10048_));
 sky130_fd_sc_hd__a21oi_4 _20311_ (.A1(_09610_),
    .A2(_09618_),
    .B1(_10046_),
    .Y(_10049_));
 sky130_fd_sc_hd__nand2_1 _20312_ (.A(_10048_),
    .B(_10045_),
    .Y(_10050_));
 sky130_fd_sc_hd__a31oi_1 _20313_ (.A1(_09610_),
    .A2(_09618_),
    .A3(_10046_),
    .B1(_05392_),
    .Y(_10051_));
 sky130_fd_sc_hd__o22ai_4 _20314_ (.A1(_05348_),
    .A2(net401),
    .B1(_10045_),
    .B2(_10048_),
    .Y(_10052_));
 sky130_fd_sc_hd__nand2_1 _20315_ (.A(_10051_),
    .B(_10050_),
    .Y(_10053_));
 sky130_fd_sc_hd__o22a_2 _20316_ (.A1(_05403_),
    .A2(_10040_),
    .B1(_10049_),
    .B2(_10052_),
    .X(_10054_));
 sky130_fd_sc_hd__o21ai_2 _20317_ (.A1(_10049_),
    .A2(_10052_),
    .B1(_10042_),
    .Y(_10055_));
 sky130_fd_sc_hd__and3_1 _20318_ (.A(_05687_),
    .B(_05709_),
    .C(_10055_),
    .X(_10056_));
 sky130_fd_sc_hd__or3_2 _20319_ (.A(_05676_),
    .B(_05698_),
    .C(_10054_),
    .X(_10057_));
 sky130_fd_sc_hd__a2bb2oi_1 _20320_ (.A1_N(_08724_),
    .A2_N(_08726_),
    .B1(_10042_),
    .B2(_10053_),
    .Y(_10059_));
 sky130_fd_sc_hd__o21ai_2 _20321_ (.A1(_08724_),
    .A2(_08726_),
    .B1(_10055_),
    .Y(_10060_));
 sky130_fd_sc_hd__o22a_1 _20322_ (.A1(_08728_),
    .A2(net195),
    .B1(_10049_),
    .B2(_10052_),
    .X(_10061_));
 sky130_fd_sc_hd__o221ai_4 _20323_ (.A1(_05403_),
    .A2(_10040_),
    .B1(_10049_),
    .B2(_10052_),
    .C1(net177),
    .Y(_10062_));
 sky130_fd_sc_hd__a21oi_2 _20324_ (.A1(_10042_),
    .A2(_10061_),
    .B1(_10059_),
    .Y(_10063_));
 sky130_fd_sc_hd__nand2_2 _20325_ (.A(_10060_),
    .B(_10062_),
    .Y(_10064_));
 sky130_fd_sc_hd__o32a_1 _20326_ (.A1(_08311_),
    .A2(_08312_),
    .A3(_09623_),
    .B1(_09643_),
    .B2(_09637_),
    .X(_10065_));
 sky130_fd_sc_hd__o22ai_2 _20327_ (.A1(net199),
    .A2(_09623_),
    .B1(_09643_),
    .B2(_09637_),
    .Y(_10066_));
 sky130_fd_sc_hd__nand2_4 _20328_ (.A(_10066_),
    .B(_10063_),
    .Y(_10067_));
 sky130_fd_sc_hd__o211ai_4 _20329_ (.A1(_09643_),
    .A2(_09637_),
    .B1(_09625_),
    .C1(_10064_),
    .Y(_10068_));
 sky130_fd_sc_hd__o221a_1 _20330_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_10063_),
    .B2(_10066_),
    .C1(_10067_),
    .X(_10070_));
 sky130_fd_sc_hd__nand3_2 _20331_ (.A(_10067_),
    .B(_10068_),
    .C(net358),
    .Y(_10071_));
 sky130_fd_sc_hd__o31a_1 _20332_ (.A1(_05676_),
    .A2(_05698_),
    .A3(_10054_),
    .B1(_10071_),
    .X(_10072_));
 sky130_fd_sc_hd__o211a_2 _20333_ (.A1(_10056_),
    .A2(_10070_),
    .B1(_06804_),
    .C1(_06826_),
    .X(_10073_));
 sky130_fd_sc_hd__or3_1 _20334_ (.A(_06793_),
    .B(_06815_),
    .C(_10072_),
    .X(_10074_));
 sky130_fd_sc_hd__a2bb2oi_4 _20335_ (.A1_N(_08307_),
    .A2_N(_08309_),
    .B1(_10057_),
    .B2(_10071_),
    .Y(_10075_));
 sky130_fd_sc_hd__o22ai_1 _20336_ (.A1(_08307_),
    .A2(_08309_),
    .B1(_10056_),
    .B2(_10070_),
    .Y(_10076_));
 sky130_fd_sc_hd__a31oi_2 _20337_ (.A1(_10067_),
    .A2(_10068_),
    .A3(net358),
    .B1(net198),
    .Y(_10077_));
 sky130_fd_sc_hd__a31o_1 _20338_ (.A1(_10067_),
    .A2(_10068_),
    .A3(net358),
    .B1(net198),
    .X(_10078_));
 sky130_fd_sc_hd__o221a_1 _20339_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_10054_),
    .B2(net358),
    .C1(_10071_),
    .X(_10079_));
 sky130_fd_sc_hd__a21oi_4 _20340_ (.A1(_10057_),
    .A2(_10077_),
    .B1(_10075_),
    .Y(_10081_));
 sky130_fd_sc_hd__nand3_1 _20341_ (.A(_08785_),
    .B(_08787_),
    .C(_08371_),
    .Y(_10082_));
 sky130_fd_sc_hd__nor3_2 _20342_ (.A(_10082_),
    .B(_09195_),
    .C(_09193_),
    .Y(_10083_));
 sky130_fd_sc_hd__nand4_1 _20343_ (.A(_09194_),
    .B(_09196_),
    .C(_08371_),
    .D(_08788_),
    .Y(_10084_));
 sky130_fd_sc_hd__a21oi_2 _20344_ (.A1(_10083_),
    .A2(_09660_),
    .B1(_09661_),
    .Y(_10085_));
 sky130_fd_sc_hd__o32ai_1 _20345_ (.A1(_07935_),
    .A2(_09651_),
    .A3(_09652_),
    .B1(_10084_),
    .B2(_09659_),
    .Y(_10086_));
 sky130_fd_sc_hd__a31oi_1 _20346_ (.A1(_09658_),
    .A2(_09660_),
    .A3(_09662_),
    .B1(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__nand2_2 _20347_ (.A(_09663_),
    .B(_10085_),
    .Y(_10088_));
 sky130_fd_sc_hd__o211ai_2 _20348_ (.A1(_07935_),
    .A2(_09655_),
    .B1(_10083_),
    .C1(_08383_),
    .Y(_10089_));
 sky130_fd_sc_hd__nand4_4 _20349_ (.A(_10083_),
    .B(_09662_),
    .C(_09660_),
    .D(_08383_),
    .Y(_10090_));
 sky130_fd_sc_hd__a2bb2oi_1 _20350_ (.A1_N(_09659_),
    .A2_N(_10089_),
    .B1(_09663_),
    .B2(_10085_),
    .Y(_10092_));
 sky130_fd_sc_hd__o2bb2ai_4 _20351_ (.A1_N(_10085_),
    .A2_N(_09663_),
    .B1(_09659_),
    .B2(_10089_),
    .Y(_10093_));
 sky130_fd_sc_hd__o211ai_1 _20352_ (.A1(_10078_),
    .A2(_10056_),
    .B1(_10076_),
    .C1(_10090_),
    .Y(_10094_));
 sky130_fd_sc_hd__nand3_4 _20353_ (.A(_10088_),
    .B(_10090_),
    .C(_10081_),
    .Y(_10095_));
 sky130_fd_sc_hd__o21ai_2 _20354_ (.A1(_10075_),
    .A2(_10079_),
    .B1(_10093_),
    .Y(_10096_));
 sky130_fd_sc_hd__o221a_1 _20355_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_10081_),
    .B2(_10092_),
    .C1(_10095_),
    .X(_10097_));
 sky130_fd_sc_hd__o221ai_2 _20356_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_10081_),
    .B2(_10092_),
    .C1(_10095_),
    .Y(_10098_));
 sky130_fd_sc_hd__o311a_2 _20357_ (.A1(_05676_),
    .A2(_05698_),
    .A3(_10054_),
    .B1(_10071_),
    .C1(_06848_),
    .X(_10099_));
 sky130_fd_sc_hd__a21oi_2 _20358_ (.A1(_10095_),
    .A2(_10096_),
    .B1(_06848_),
    .Y(_10100_));
 sky130_fd_sc_hd__a31oi_4 _20359_ (.A1(_10096_),
    .A2(net357),
    .A3(_10095_),
    .B1(_10073_),
    .Y(_10101_));
 sky130_fd_sc_hd__a21oi_2 _20360_ (.A1(_09678_),
    .A2(_09681_),
    .B1(_09672_),
    .Y(_10103_));
 sky130_fd_sc_hd__o32ai_4 _20361_ (.A1(_07564_),
    .A2(_09667_),
    .A3(_09668_),
    .B1(_09679_),
    .B2(_09680_),
    .Y(_10104_));
 sky130_fd_sc_hd__a2bb2oi_1 _20362_ (.A1_N(_07928_),
    .A2_N(_07930_),
    .B1(_09673_),
    .B2(_09683_),
    .Y(_10105_));
 sky130_fd_sc_hd__a31oi_2 _20363_ (.A1(_09683_),
    .A2(_07935_),
    .A3(_09673_),
    .B1(_07724_),
    .Y(_10106_));
 sky130_fd_sc_hd__o22ai_2 _20364_ (.A1(_07691_),
    .A2(net371),
    .B1(_07936_),
    .B2(_10104_),
    .Y(_10107_));
 sky130_fd_sc_hd__o221ai_4 _20365_ (.A1(_10073_),
    .A2(_10097_),
    .B1(_10103_),
    .B2(_07935_),
    .C1(_10106_),
    .Y(_10108_));
 sky130_fd_sc_hd__o22ai_4 _20366_ (.A1(_10099_),
    .A2(_10100_),
    .B1(_10105_),
    .B2(_10107_),
    .Y(_10109_));
 sky130_fd_sc_hd__or4_2 _20367_ (.A(net374),
    .B(_07702_),
    .C(_10099_),
    .D(_10100_),
    .X(_10110_));
 sky130_fd_sc_hd__o211a_1 _20368_ (.A1(net357),
    .A2(_10072_),
    .B1(_07935_),
    .C1(_10098_),
    .X(_10111_));
 sky130_fd_sc_hd__a311o_1 _20369_ (.A1(_10096_),
    .A2(net357),
    .A3(_10095_),
    .B1(_07936_),
    .C1(_10073_),
    .X(_10112_));
 sky130_fd_sc_hd__a21oi_1 _20370_ (.A1(_10074_),
    .A2(_10098_),
    .B1(_07935_),
    .Y(_10114_));
 sky130_fd_sc_hd__o21ai_1 _20371_ (.A1(_10073_),
    .A2(_10097_),
    .B1(_07936_),
    .Y(_10115_));
 sky130_fd_sc_hd__nand3_2 _20372_ (.A(_10104_),
    .B(_10112_),
    .C(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__o21ai_2 _20373_ (.A1(_10111_),
    .A2(_10114_),
    .B1(_10103_),
    .Y(_10117_));
 sky130_fd_sc_hd__nand3_4 _20374_ (.A(_10117_),
    .B(net354),
    .C(_10116_),
    .Y(_10118_));
 sky130_fd_sc_hd__o31a_1 _20375_ (.A1(net354),
    .A2(_10099_),
    .A3(_10100_),
    .B1(_10118_),
    .X(_10119_));
 sky130_fd_sc_hd__a2bb2oi_4 _20376_ (.A1_N(_07555_),
    .A2_N(net218),
    .B1(_10110_),
    .B2(_10118_),
    .Y(_10120_));
 sky130_fd_sc_hd__o211ai_4 _20377_ (.A1(_07555_),
    .A2(net218),
    .B1(_10108_),
    .C1(_10109_),
    .Y(_10121_));
 sky130_fd_sc_hd__a31oi_1 _20378_ (.A1(_10117_),
    .A2(net354),
    .A3(_10116_),
    .B1(net202),
    .Y(_10122_));
 sky130_fd_sc_hd__o311a_1 _20379_ (.A1(net354),
    .A2(_10099_),
    .A3(_10100_),
    .B1(_07564_),
    .C1(_10118_),
    .X(_10123_));
 sky130_fd_sc_hd__o211ai_4 _20380_ (.A1(net354),
    .A2(_10101_),
    .B1(_07564_),
    .C1(_10118_),
    .Y(_10125_));
 sky130_fd_sc_hd__a21oi_1 _20381_ (.A1(_10110_),
    .A2(_10122_),
    .B1(_10120_),
    .Y(_10126_));
 sky130_fd_sc_hd__o211ai_4 _20382_ (.A1(_09693_),
    .A2(_09239_),
    .B1(_09229_),
    .C1(_09690_),
    .Y(_10127_));
 sky130_fd_sc_hd__o21ai_1 _20383_ (.A1(net222),
    .A2(_09688_),
    .B1(_10127_),
    .Y(_10128_));
 sky130_fd_sc_hd__o21ai_4 _20384_ (.A1(_10120_),
    .A2(_10123_),
    .B1(_10128_),
    .Y(_10129_));
 sky130_fd_sc_hd__nand4_4 _20385_ (.A(_09692_),
    .B(_10121_),
    .C(_10125_),
    .D(_10127_),
    .Y(_10130_));
 sky130_fd_sc_hd__and3_2 _20386_ (.A(_08732_),
    .B(_10108_),
    .C(_10109_),
    .X(_10131_));
 sky130_fd_sc_hd__inv_2 _20387_ (.A(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__nand3_1 _20388_ (.A(_10129_),
    .B(_10130_),
    .C(net338),
    .Y(_10133_));
 sky130_fd_sc_hd__a31o_1 _20389_ (.A1(_10129_),
    .A2(_10130_),
    .A3(net338),
    .B1(_10131_),
    .X(_10134_));
 sky130_fd_sc_hd__a31oi_4 _20390_ (.A1(_10129_),
    .A2(_10130_),
    .A3(net338),
    .B1(_10131_),
    .Y(_10136_));
 sky130_fd_sc_hd__a2bb2oi_2 _20391_ (.A1_N(_07242_),
    .A2_N(_07243_),
    .B1(_10132_),
    .B2(_10133_),
    .Y(_10137_));
 sky130_fd_sc_hd__a2bb2o_1 _20392_ (.A1_N(_07242_),
    .A2_N(_07243_),
    .B1(_10132_),
    .B2(_10133_),
    .X(_10138_));
 sky130_fd_sc_hd__a311oi_4 _20393_ (.A1(_10129_),
    .A2(_10130_),
    .A3(net338),
    .B1(_10131_),
    .C1(net222),
    .Y(_10139_));
 sky130_fd_sc_hd__a311o_1 _20394_ (.A1(_10129_),
    .A2(_10130_),
    .A3(net338),
    .B1(_10131_),
    .C1(net222),
    .X(_10140_));
 sky130_fd_sc_hd__o2bb2ai_1 _20395_ (.A1_N(_09715_),
    .A2_N(_09717_),
    .B1(net227),
    .B2(_09704_),
    .Y(_10141_));
 sky130_fd_sc_hd__o211ai_2 _20396_ (.A1(net225),
    .A2(_09703_),
    .B1(_09715_),
    .C1(_09717_),
    .Y(_10142_));
 sky130_fd_sc_hd__o221ai_4 _20397_ (.A1(_09704_),
    .A2(net227),
    .B1(_10139_),
    .B2(_10137_),
    .C1(_09725_),
    .Y(_10143_));
 sky130_fd_sc_hd__o2111ai_4 _20398_ (.A1(_09703_),
    .A2(net225),
    .B1(_10140_),
    .C1(_10138_),
    .D1(_10141_),
    .Y(_10144_));
 sky130_fd_sc_hd__nand3_4 _20399_ (.A(_10144_),
    .B(net335),
    .C(_10143_),
    .Y(_10145_));
 sky130_fd_sc_hd__or3_2 _20400_ (.A(net351),
    .B(_09807_),
    .C(_10136_),
    .X(_10147_));
 sky130_fd_sc_hd__o21ai_4 _20401_ (.A1(net335),
    .A2(_10136_),
    .B1(_10145_),
    .Y(_10148_));
 sky130_fd_sc_hd__inv_2 _20402_ (.A(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__o311a_1 _20403_ (.A1(net351),
    .A2(_10136_),
    .A3(_09807_),
    .B1(_11079_),
    .C1(_10145_),
    .X(_10150_));
 sky130_fd_sc_hd__a22oi_4 _20404_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_10145_),
    .B2(_10147_),
    .Y(_10151_));
 sky130_fd_sc_hd__a21o_1 _20405_ (.A1(_10145_),
    .A2(_10147_),
    .B1(net227),
    .X(_10152_));
 sky130_fd_sc_hd__o221a_1 _20406_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_10136_),
    .B2(net335),
    .C1(_10145_),
    .X(_10153_));
 sky130_fd_sc_hd__o221ai_4 _20407_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_10136_),
    .B2(net336),
    .C1(_10145_),
    .Y(_10154_));
 sky130_fd_sc_hd__nor2_1 _20408_ (.A(_10151_),
    .B(_10153_),
    .Y(_10155_));
 sky130_fd_sc_hd__nand2_1 _20409_ (.A(_10152_),
    .B(_10154_),
    .Y(_10156_));
 sky130_fd_sc_hd__and3_1 _20410_ (.A(_08462_),
    .B(_08860_),
    .C(_08861_),
    .X(_10158_));
 sky130_fd_sc_hd__o211a_1 _20411_ (.A1(_09252_),
    .A2(_09273_),
    .B1(_10158_),
    .C1(_09271_),
    .X(_10159_));
 sky130_fd_sc_hd__nand3_1 _20412_ (.A(_09732_),
    .B(_10158_),
    .C(_09276_),
    .Y(_10160_));
 sky130_fd_sc_hd__nand4_2 _20413_ (.A(_09732_),
    .B(_09733_),
    .C(_10158_),
    .D(_09276_),
    .Y(_10161_));
 sky130_fd_sc_hd__nand4_4 _20414_ (.A(_10159_),
    .B(_09733_),
    .C(_09732_),
    .D(_08454_),
    .Y(_10162_));
 sky130_fd_sc_hd__o211a_1 _20415_ (.A1(_09736_),
    .A2(_09731_),
    .B1(_09733_),
    .C1(_10160_),
    .X(_10163_));
 sky130_fd_sc_hd__o211ai_4 _20416_ (.A1(_09736_),
    .A2(_09731_),
    .B1(_09733_),
    .C1(_10160_),
    .Y(_10164_));
 sky130_fd_sc_hd__o21ai_2 _20417_ (.A1(_08455_),
    .A2(_10161_),
    .B1(_10164_),
    .Y(_10165_));
 sky130_fd_sc_hd__a21oi_2 _20418_ (.A1(_10162_),
    .A2(_10164_),
    .B1(_10156_),
    .Y(_10166_));
 sky130_fd_sc_hd__nand2_1 _20419_ (.A(_10165_),
    .B(_10155_),
    .Y(_10167_));
 sky130_fd_sc_hd__o211ai_2 _20420_ (.A1(_10151_),
    .A2(_10153_),
    .B1(_10162_),
    .C1(_10164_),
    .Y(_10169_));
 sky130_fd_sc_hd__o21ai_2 _20421_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__a211o_1 _20422_ (.A1(_10145_),
    .A2(_10147_),
    .B1(_11046_),
    .C1(_11057_),
    .X(_10171_));
 sky130_fd_sc_hd__inv_2 _20423_ (.A(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__nand4_4 _20424_ (.A(_10152_),
    .B(_10154_),
    .C(_10162_),
    .D(_10164_),
    .Y(_10173_));
 sky130_fd_sc_hd__o21ai_2 _20425_ (.A1(_10151_),
    .A2(_10153_),
    .B1(_10165_),
    .Y(_10174_));
 sky130_fd_sc_hd__nand3_1 _20426_ (.A(_10174_),
    .B(net333),
    .C(_10173_),
    .Y(_10175_));
 sky130_fd_sc_hd__o221a_2 _20427_ (.A1(net333),
    .A2(_10148_),
    .B1(_10166_),
    .B2(_10170_),
    .C1(_12703_),
    .X(_10176_));
 sky130_fd_sc_hd__a311o_2 _20428_ (.A1(_10167_),
    .A2(_10169_),
    .A3(net333),
    .B1(net311),
    .C1(_10150_),
    .X(_10177_));
 sky130_fd_sc_hd__a311oi_4 _20429_ (.A1(_10174_),
    .A2(net333),
    .A3(_10173_),
    .B1(net232),
    .C1(_10172_),
    .Y(_10178_));
 sky130_fd_sc_hd__nand3_4 _20430_ (.A(_10175_),
    .B(net234),
    .C(_10171_),
    .Y(_10180_));
 sky130_fd_sc_hd__a311oi_1 _20431_ (.A1(_10167_),
    .A2(_10169_),
    .A3(net333),
    .B1(net234),
    .C1(_10150_),
    .Y(_10181_));
 sky130_fd_sc_hd__o221ai_4 _20432_ (.A1(net333),
    .A2(_10148_),
    .B1(_10166_),
    .B2(_10170_),
    .C1(net232),
    .Y(_10182_));
 sky130_fd_sc_hd__a211oi_1 _20433_ (.A1(_09293_),
    .A2(_09290_),
    .B1(_09287_),
    .C1(_09747_),
    .Y(_10183_));
 sky130_fd_sc_hd__a22oi_2 _20434_ (.A1(_09729_),
    .A2(_09743_),
    .B1(_09740_),
    .B2(_09748_),
    .Y(_10184_));
 sky130_fd_sc_hd__o22ai_2 _20435_ (.A1(_09728_),
    .A2(_09744_),
    .B1(_09747_),
    .B2(_09742_),
    .Y(_10185_));
 sky130_fd_sc_hd__o2bb2ai_2 _20436_ (.A1_N(_10180_),
    .A2_N(_10182_),
    .B1(_10183_),
    .B2(_09745_),
    .Y(_10186_));
 sky130_fd_sc_hd__nand3_4 _20437_ (.A(_10184_),
    .B(_10182_),
    .C(_10180_),
    .Y(_10187_));
 sky130_fd_sc_hd__nand3_2 _20438_ (.A(_10186_),
    .B(_10187_),
    .C(net312),
    .Y(_10188_));
 sky130_fd_sc_hd__a31o_2 _20439_ (.A1(_10186_),
    .A2(_10187_),
    .A3(net311),
    .B1(_10176_),
    .X(_10189_));
 sky130_fd_sc_hd__nand2_1 _20440_ (.A(_09758_),
    .B(_09766_),
    .Y(_10191_));
 sky130_fd_sc_hd__o2bb2ai_1 _20441_ (.A1_N(_09314_),
    .A2_N(_09764_),
    .B1(_09756_),
    .B2(net253),
    .Y(_10192_));
 sky130_fd_sc_hd__o21bai_1 _20442_ (.A1(_09760_),
    .A2(_09766_),
    .B1_N(_09757_),
    .Y(_10193_));
 sky130_fd_sc_hd__a311oi_4 _20443_ (.A1(_10186_),
    .A2(_10187_),
    .A3(net311),
    .B1(net251),
    .C1(_10176_),
    .Y(_10194_));
 sky130_fd_sc_hd__o211ai_4 _20444_ (.A1(_06309_),
    .A2(_06312_),
    .B1(_10177_),
    .C1(_10188_),
    .Y(_10195_));
 sky130_fd_sc_hd__a21oi_2 _20445_ (.A1(_10177_),
    .A2(_10188_),
    .B1(_06314_),
    .Y(_10196_));
 sky130_fd_sc_hd__a22o_1 _20446_ (.A1(_06306_),
    .A2(_06308_),
    .B1(_10177_),
    .B2(_10188_),
    .X(_10197_));
 sky130_fd_sc_hd__o2111ai_4 _20447_ (.A1(_09760_),
    .A2(_09766_),
    .B1(_10195_),
    .C1(_10197_),
    .D1(_09758_),
    .Y(_10198_));
 sky130_fd_sc_hd__o21ai_1 _20448_ (.A1(_10194_),
    .A2(_10196_),
    .B1(_10193_),
    .Y(_10199_));
 sky130_fd_sc_hd__nand3_4 _20449_ (.A(_10198_),
    .B(_10199_),
    .C(net308),
    .Y(_10200_));
 sky130_fd_sc_hd__a211o_1 _20450_ (.A1(_10177_),
    .A2(_10188_),
    .B1(_00011_),
    .C1(net323),
    .X(_10202_));
 sky130_fd_sc_hd__o2111ai_4 _20451_ (.A1(net253),
    .A2(_09756_),
    .B1(_10191_),
    .C1(_10195_),
    .D1(_10197_),
    .Y(_10203_));
 sky130_fd_sc_hd__o2bb2ai_1 _20452_ (.A1_N(_09761_),
    .A2_N(_10191_),
    .B1(_10194_),
    .B2(_10196_),
    .Y(_10204_));
 sky130_fd_sc_hd__o211ai_4 _20453_ (.A1(_00011_),
    .A2(net323),
    .B1(_10203_),
    .C1(_10204_),
    .Y(_10205_));
 sky130_fd_sc_hd__o21ai_4 _20454_ (.A1(net307),
    .A2(_10189_),
    .B1(_10200_),
    .Y(_10206_));
 sky130_fd_sc_hd__o211ai_4 _20455_ (.A1(_10189_),
    .A2(net307),
    .B1(net253),
    .C1(_10200_),
    .Y(_10207_));
 sky130_fd_sc_hd__and3_2 _20456_ (.A(_10205_),
    .B(net254),
    .C(_10202_),
    .X(_10208_));
 sky130_fd_sc_hd__o211ai_4 _20457_ (.A1(net286),
    .A2(_06012_),
    .B1(_10202_),
    .C1(_10205_),
    .Y(_10209_));
 sky130_fd_sc_hd__nand2_1 _20458_ (.A(_10207_),
    .B(_10209_),
    .Y(_10210_));
 sky130_fd_sc_hd__a21o_1 _20459_ (.A1(_09783_),
    .A2(_09787_),
    .B1(_09777_),
    .X(_10211_));
 sky130_fd_sc_hd__nand3_2 _20460_ (.A(_09779_),
    .B(_09783_),
    .C(_09787_),
    .Y(_10213_));
 sky130_fd_sc_hd__a31oi_2 _20461_ (.A1(_09779_),
    .A2(_09783_),
    .A3(_09787_),
    .B1(_09777_),
    .Y(_10214_));
 sky130_fd_sc_hd__a22oi_4 _20462_ (.A1(_10207_),
    .A2(_10209_),
    .B1(_10211_),
    .B2(_09779_),
    .Y(_10215_));
 sky130_fd_sc_hd__o22ai_4 _20463_ (.A1(_01940_),
    .A2(_01951_),
    .B1(_10210_),
    .B2(_10214_),
    .Y(_10216_));
 sky130_fd_sc_hd__o22ai_4 _20464_ (.A1(net279),
    .A2(_10206_),
    .B1(_10215_),
    .B2(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__o21a_1 _20465_ (.A1(_05760_),
    .A2(net290),
    .B1(_10217_),
    .X(_10218_));
 sky130_fd_sc_hd__o21ai_4 _20466_ (.A1(_05760_),
    .A2(net290),
    .B1(_10217_),
    .Y(_10219_));
 sky130_fd_sc_hd__o221ai_4 _20467_ (.A1(net279),
    .A2(_10206_),
    .B1(_10215_),
    .B2(_10216_),
    .C1(net262),
    .Y(_10220_));
 sky130_fd_sc_hd__and3_1 _20468_ (.A(_08935_),
    .B(_08937_),
    .C(_08528_),
    .X(_10221_));
 sky130_fd_sc_hd__nand3_1 _20469_ (.A(_09802_),
    .B(_10221_),
    .C(_09350_),
    .Y(_10222_));
 sky130_fd_sc_hd__o211ai_4 _20470_ (.A1(_09806_),
    .A2(_09801_),
    .B1(_09803_),
    .C1(_10222_),
    .Y(_10224_));
 sky130_fd_sc_hd__and4_1 _20471_ (.A(_10221_),
    .B(_09349_),
    .C(_09347_),
    .D(_08536_),
    .X(_10225_));
 sky130_fd_sc_hd__nand3_4 _20472_ (.A(_10225_),
    .B(_09803_),
    .C(_09802_),
    .Y(_10226_));
 sky130_fd_sc_hd__and2_2 _20473_ (.A(_10224_),
    .B(_10226_),
    .X(_10227_));
 sky130_fd_sc_hd__o211ai_4 _20474_ (.A1(net261),
    .A2(_10217_),
    .B1(_10224_),
    .C1(_10226_),
    .Y(_10228_));
 sky130_fd_sc_hd__o2111ai_4 _20475_ (.A1(net261),
    .A2(_10217_),
    .B1(_10219_),
    .C1(_10224_),
    .D1(_10226_),
    .Y(_10229_));
 sky130_fd_sc_hd__a22o_2 _20476_ (.A1(_10219_),
    .A2(_10220_),
    .B1(_10224_),
    .B2(_10226_),
    .X(_10230_));
 sky130_fd_sc_hd__nand3_1 _20477_ (.A(_10230_),
    .B(net276),
    .C(_10229_),
    .Y(_10231_));
 sky130_fd_sc_hd__o21a_2 _20478_ (.A1(_03986_),
    .A2(_03997_),
    .B1(_10217_),
    .X(_10232_));
 sky130_fd_sc_hd__o21ai_1 _20479_ (.A1(_03986_),
    .A2(_03997_),
    .B1(_10217_),
    .Y(_10233_));
 sky130_fd_sc_hd__a31oi_4 _20480_ (.A1(_10230_),
    .A2(net276),
    .A3(_10229_),
    .B1(_10232_),
    .Y(_10235_));
 sky130_fd_sc_hd__a2bb2o_2 _20481_ (.A1_N(_05228_),
    .A2_N(_05230_),
    .B1(_10231_),
    .B2(_10233_),
    .X(_10236_));
 sky130_fd_sc_hd__inv_2 _20482_ (.A(_10236_),
    .Y(_10237_));
 sky130_fd_sc_hd__a31o_1 _20483_ (.A1(_10230_),
    .A2(net276),
    .A3(_10229_),
    .B1(net291),
    .X(_10238_));
 sky130_fd_sc_hd__a311oi_4 _20484_ (.A1(_10230_),
    .A2(net276),
    .A3(_10229_),
    .B1(_10232_),
    .C1(net291),
    .Y(_10239_));
 sky130_fd_sc_hd__nand3_1 _20485_ (.A(_10231_),
    .B(_10233_),
    .C(net267),
    .Y(_10240_));
 sky130_fd_sc_hd__a21oi_1 _20486_ (.A1(_10231_),
    .A2(_10233_),
    .B1(net267),
    .Y(_10241_));
 sky130_fd_sc_hd__a22o_2 _20487_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_10231_),
    .B2(_10233_),
    .X(_10242_));
 sky130_fd_sc_hd__o2bb2a_1 _20488_ (.A1_N(_09821_),
    .A2_N(_09800_),
    .B1(_09820_),
    .B2(_09824_),
    .X(_10243_));
 sky130_fd_sc_hd__a21oi_2 _20489_ (.A1(_09823_),
    .A2(_09820_),
    .B1(_09824_),
    .Y(_10244_));
 sky130_fd_sc_hd__o21a_1 _20490_ (.A1(_10239_),
    .A2(_10241_),
    .B1(_10244_),
    .X(_10246_));
 sky130_fd_sc_hd__o21ai_2 _20491_ (.A1(_10239_),
    .A2(_10241_),
    .B1(_10244_),
    .Y(_10247_));
 sky130_fd_sc_hd__o21ai_2 _20492_ (.A1(net267),
    .A2(_10235_),
    .B1(_10243_),
    .Y(_10248_));
 sky130_fd_sc_hd__o211ai_2 _20493_ (.A1(_10232_),
    .A2(_10238_),
    .B1(_10243_),
    .C1(_10242_),
    .Y(_10249_));
 sky130_fd_sc_hd__o21ai_2 _20494_ (.A1(_10239_),
    .A2(_10248_),
    .B1(net273),
    .Y(_10250_));
 sky130_fd_sc_hd__o211ai_4 _20495_ (.A1(_10239_),
    .A2(_10248_),
    .B1(net273),
    .C1(_10247_),
    .Y(_10251_));
 sky130_fd_sc_hd__o22ai_4 _20496_ (.A1(net273),
    .A2(_10235_),
    .B1(_10246_),
    .B2(_10250_),
    .Y(_10252_));
 sky130_fd_sc_hd__o221a_1 _20497_ (.A1(net273),
    .A2(_10235_),
    .B1(_10246_),
    .B2(_10250_),
    .C1(_05486_),
    .X(_10253_));
 sky130_fd_sc_hd__o2bb2a_1 _20498_ (.A1_N(net298),
    .A2_N(_09834_),
    .B1(_09839_),
    .B2(_09376_),
    .X(_10254_));
 sky130_fd_sc_hd__o211a_1 _20499_ (.A1(_02148_),
    .A2(_09373_),
    .B1(_09838_),
    .C1(_09841_),
    .X(_10255_));
 sky130_fd_sc_hd__a31o_1 _20500_ (.A1(_09377_),
    .A2(_09838_),
    .A3(_09841_),
    .B1(_09835_),
    .X(_10257_));
 sky130_fd_sc_hd__a311oi_4 _20501_ (.A1(_10247_),
    .A2(_10249_),
    .A3(net273),
    .B1(net294),
    .C1(_10237_),
    .Y(_10258_));
 sky130_fd_sc_hd__o211ai_4 _20502_ (.A1(net273),
    .A2(_10235_),
    .B1(net295),
    .C1(_10251_),
    .Y(_10259_));
 sky130_fd_sc_hd__a2bb2oi_2 _20503_ (.A1_N(net318),
    .A2_N(_05244_),
    .B1(_10236_),
    .B2(_10251_),
    .Y(_10260_));
 sky130_fd_sc_hd__a22o_1 _20504_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_10236_),
    .B2(_10251_),
    .X(_10261_));
 sky130_fd_sc_hd__o211ai_2 _20505_ (.A1(_09837_),
    .A2(_10254_),
    .B1(_10259_),
    .C1(_10261_),
    .Y(_10262_));
 sky130_fd_sc_hd__o22ai_2 _20506_ (.A1(_09835_),
    .A2(_10255_),
    .B1(_10258_),
    .B2(_10260_),
    .Y(_10263_));
 sky130_fd_sc_hd__nand3_1 _20507_ (.A(_10262_),
    .B(_10263_),
    .C(net246),
    .Y(_10264_));
 sky130_fd_sc_hd__a211o_1 _20508_ (.A1(_10236_),
    .A2(_10251_),
    .B1(_05481_),
    .C1(_05483_),
    .X(_10265_));
 sky130_fd_sc_hd__o211ai_1 _20509_ (.A1(_09835_),
    .A2(_10255_),
    .B1(_10259_),
    .C1(_10261_),
    .Y(_10266_));
 sky130_fd_sc_hd__o22ai_1 _20510_ (.A1(_09837_),
    .A2(_10254_),
    .B1(_10258_),
    .B2(_10260_),
    .Y(_10268_));
 sky130_fd_sc_hd__nand3_1 _20511_ (.A(_10266_),
    .B(_10268_),
    .C(net246),
    .Y(_10269_));
 sky130_fd_sc_hd__a31o_2 _20512_ (.A1(_10262_),
    .A2(_10263_),
    .A3(net246),
    .B1(_10253_),
    .X(_10270_));
 sky130_fd_sc_hd__nand2_1 _20513_ (.A(_05754_),
    .B(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__o211ai_4 _20514_ (.A1(_10252_),
    .A2(net246),
    .B1(net298),
    .C1(_10264_),
    .Y(_10272_));
 sky130_fd_sc_hd__and3_1 _20515_ (.A(_10269_),
    .B(net299),
    .C(_10265_),
    .X(_10273_));
 sky130_fd_sc_hd__nand3_4 _20516_ (.A(_10269_),
    .B(net299),
    .C(_10265_),
    .Y(_10274_));
 sky130_fd_sc_hd__a21oi_1 _20517_ (.A1(_02148_),
    .A2(_09847_),
    .B1(_09854_),
    .Y(_10275_));
 sky130_fd_sc_hd__o21ai_2 _20518_ (.A1(_09855_),
    .A2(_09852_),
    .B1(_09850_),
    .Y(_10276_));
 sky130_fd_sc_hd__o2111ai_1 _20519_ (.A1(_09855_),
    .A2(_09852_),
    .B1(_09850_),
    .C1(_10274_),
    .D1(_10272_),
    .Y(_10277_));
 sky130_fd_sc_hd__a22o_1 _20520_ (.A1(_09850_),
    .A2(_09856_),
    .B1(_10272_),
    .B2(_10274_),
    .X(_10279_));
 sky130_fd_sc_hd__o211ai_2 _20521_ (.A1(net266),
    .A2(_05751_),
    .B1(_10277_),
    .C1(_10279_),
    .Y(_10280_));
 sky130_fd_sc_hd__o211a_1 _20522_ (.A1(_10252_),
    .A2(net246),
    .B1(_05754_),
    .C1(_10264_),
    .X(_10281_));
 sky130_fd_sc_hd__a311o_1 _20523_ (.A1(_10262_),
    .A2(_10263_),
    .A3(net246),
    .B1(net242),
    .C1(_10253_),
    .X(_10282_));
 sky130_fd_sc_hd__a21oi_2 _20524_ (.A1(_10272_),
    .A2(_10274_),
    .B1(_10276_),
    .Y(_10283_));
 sky130_fd_sc_hd__o2bb2ai_1 _20525_ (.A1_N(_10272_),
    .A2_N(_10274_),
    .B1(_10275_),
    .B2(_09852_),
    .Y(_10284_));
 sky130_fd_sc_hd__nand3_1 _20526_ (.A(_10272_),
    .B(_10274_),
    .C(_10276_),
    .Y(_10285_));
 sky130_fd_sc_hd__a31o_1 _20527_ (.A1(_10272_),
    .A2(_10274_),
    .A3(_10276_),
    .B1(_05754_),
    .X(_10286_));
 sky130_fd_sc_hd__nand3_1 _20528_ (.A(_10284_),
    .B(_10285_),
    .C(net242),
    .Y(_10287_));
 sky130_fd_sc_hd__a311o_2 _20529_ (.A1(_10284_),
    .A2(_10285_),
    .A3(net242),
    .B1(net240),
    .C1(_10281_),
    .X(_10288_));
 sky130_fd_sc_hd__a2bb2oi_2 _20530_ (.A1_N(_02049_),
    .A2_N(net343),
    .B1(_10282_),
    .B2(_10287_),
    .Y(_10290_));
 sky130_fd_sc_hd__o211ai_4 _20531_ (.A1(_02049_),
    .A2(net343),
    .B1(_10271_),
    .C1(_10280_),
    .Y(_10291_));
 sky130_fd_sc_hd__a31o_1 _20532_ (.A1(_10284_),
    .A2(_10285_),
    .A3(net242),
    .B1(_02148_),
    .X(_10292_));
 sky130_fd_sc_hd__o221a_1 _20533_ (.A1(net242),
    .A2(_10270_),
    .B1(_10283_),
    .B2(_10286_),
    .C1(_02137_),
    .X(_10293_));
 sky130_fd_sc_hd__o221ai_4 _20534_ (.A1(net242),
    .A2(_10270_),
    .B1(_10283_),
    .B2(_10286_),
    .C1(_02137_),
    .Y(_10294_));
 sky130_fd_sc_hd__nand4_2 _20535_ (.A(_08602_),
    .B(_08604_),
    .C(_09000_),
    .D(_09002_),
    .Y(_10295_));
 sky130_fd_sc_hd__a21oi_2 _20536_ (.A1(net326),
    .A2(_09408_),
    .B1(_10295_),
    .Y(_10296_));
 sky130_fd_sc_hd__a211oi_1 _20537_ (.A1(_09394_),
    .A2(_09415_),
    .B1(_10295_),
    .C1(_09418_),
    .Y(_10297_));
 sky130_fd_sc_hd__nand3_1 _20538_ (.A(_10296_),
    .B(_09871_),
    .C(_09417_),
    .Y(_10298_));
 sky130_fd_sc_hd__a31oi_2 _20539_ (.A1(_10296_),
    .A2(_09871_),
    .A3(_09417_),
    .B1(_09872_),
    .Y(_10299_));
 sky130_fd_sc_hd__o211a_1 _20540_ (.A1(_09878_),
    .A2(_09870_),
    .B1(_09874_),
    .C1(_10298_),
    .X(_10301_));
 sky130_fd_sc_hd__o211ai_4 _20541_ (.A1(_09878_),
    .A2(_09870_),
    .B1(_09874_),
    .C1(_10298_),
    .Y(_10302_));
 sky130_fd_sc_hd__nand4_4 _20542_ (.A(_10296_),
    .B(_09874_),
    .C(_09871_),
    .D(_09417_),
    .Y(_10303_));
 sky130_fd_sc_hd__and4_1 _20543_ (.A(_09871_),
    .B(_10297_),
    .C(_09874_),
    .D(_08606_),
    .X(_10304_));
 sky130_fd_sc_hd__nand4_1 _20544_ (.A(_09871_),
    .B(_10297_),
    .C(_09874_),
    .D(_08606_),
    .Y(_10305_));
 sky130_fd_sc_hd__a2bb2oi_4 _20545_ (.A1_N(_08607_),
    .A2_N(_10303_),
    .B1(_09882_),
    .B2(_10299_),
    .Y(_10306_));
 sky130_fd_sc_hd__o21ai_4 _20546_ (.A1(_08607_),
    .A2(_10303_),
    .B1(_10302_),
    .Y(_10307_));
 sky130_fd_sc_hd__o211ai_2 _20547_ (.A1(_10292_),
    .A2(_10281_),
    .B1(_10291_),
    .C1(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__o21ai_1 _20548_ (.A1(_10290_),
    .A2(_10293_),
    .B1(_10306_),
    .Y(_10309_));
 sky130_fd_sc_hd__o211ai_4 _20549_ (.A1(net259),
    .A2(net257),
    .B1(_10308_),
    .C1(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__and3_1 _20550_ (.A(_10280_),
    .B(_05995_),
    .C(_10271_),
    .X(_10312_));
 sky130_fd_sc_hd__a211o_2 _20551_ (.A1(_10282_),
    .A2(_10287_),
    .B1(net259),
    .C1(_05992_),
    .X(_10313_));
 sky130_fd_sc_hd__o2bb2ai_2 _20552_ (.A1_N(_10291_),
    .A2_N(_10294_),
    .B1(_10301_),
    .B2(_10304_),
    .Y(_10314_));
 sky130_fd_sc_hd__o211ai_4 _20553_ (.A1(_08607_),
    .A2(_10303_),
    .B1(_10302_),
    .C1(_10294_),
    .Y(_10315_));
 sky130_fd_sc_hd__o2111ai_2 _20554_ (.A1(_08607_),
    .A2(_10303_),
    .B1(_10302_),
    .C1(_10294_),
    .D1(_10291_),
    .Y(_10316_));
 sky130_fd_sc_hd__o221ai_4 _20555_ (.A1(net259),
    .A2(net257),
    .B1(_10290_),
    .B2(_10315_),
    .C1(_10314_),
    .Y(_10317_));
 sky130_fd_sc_hd__a31o_1 _20556_ (.A1(net240),
    .A2(_10314_),
    .A3(_10316_),
    .B1(_10312_),
    .X(_10318_));
 sky130_fd_sc_hd__inv_2 _20557_ (.A(_10318_),
    .Y(_10319_));
 sky130_fd_sc_hd__and3_1 _20558_ (.A(_06294_),
    .B(_10288_),
    .C(_10310_),
    .X(_10320_));
 sky130_fd_sc_hd__a22o_1 _20559_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_10313_),
    .B2(_10317_),
    .X(_10321_));
 sky130_fd_sc_hd__a311oi_2 _20560_ (.A1(net240),
    .A2(_10314_),
    .A3(_10316_),
    .B1(_10312_),
    .C1(_00251_),
    .Y(_10323_));
 sky130_fd_sc_hd__nand3_4 _20561_ (.A(_10317_),
    .B(_00240_),
    .C(_10313_),
    .Y(_10324_));
 sky130_fd_sc_hd__a2bb2oi_4 _20562_ (.A1_N(_00174_),
    .A2_N(net344),
    .B1(_10313_),
    .B2(_10317_),
    .Y(_10325_));
 sky130_fd_sc_hd__o211ai_4 _20563_ (.A1(_00174_),
    .A2(net344),
    .B1(_10288_),
    .C1(_10310_),
    .Y(_10326_));
 sky130_fd_sc_hd__o311a_1 _20564_ (.A1(_09018_),
    .A2(_09432_),
    .A3(_09435_),
    .B1(_09892_),
    .C1(_09431_),
    .X(_10327_));
 sky130_fd_sc_hd__o31a_1 _20565_ (.A1(_09430_),
    .A2(_09888_),
    .A3(_09891_),
    .B1(_09890_),
    .X(_10328_));
 sky130_fd_sc_hd__o31a_1 _20566_ (.A1(_09432_),
    .A2(_09887_),
    .A3(_09889_),
    .B1(_09892_),
    .X(_10329_));
 sky130_fd_sc_hd__a21oi_1 _20567_ (.A1(_10324_),
    .A2(_10326_),
    .B1(_10328_),
    .Y(_10330_));
 sky130_fd_sc_hd__o2bb2ai_2 _20568_ (.A1_N(_10324_),
    .A2_N(_10326_),
    .B1(_10327_),
    .B2(_09889_),
    .Y(_10331_));
 sky130_fd_sc_hd__nand3_2 _20569_ (.A(_10324_),
    .B(_10326_),
    .C(_10328_),
    .Y(_10332_));
 sky130_fd_sc_hd__a31o_1 _20570_ (.A1(_10324_),
    .A2(_10326_),
    .A3(_10328_),
    .B1(_06294_),
    .X(_10334_));
 sky130_fd_sc_hd__nand3_1 _20571_ (.A(_10331_),
    .B(_10332_),
    .C(net212),
    .Y(_10335_));
 sky130_fd_sc_hd__o22ai_4 _20572_ (.A1(net212),
    .A2(_10319_),
    .B1(_10330_),
    .B2(_10334_),
    .Y(_10336_));
 sky130_fd_sc_hd__o221a_1 _20573_ (.A1(_09450_),
    .A2(_09453_),
    .B1(_11298_),
    .B2(_09902_),
    .C1(_09449_),
    .X(_10337_));
 sky130_fd_sc_hd__o311a_1 _20574_ (.A1(_09034_),
    .A2(_09448_),
    .A3(_09452_),
    .B1(_09906_),
    .C1(_09451_),
    .X(_10338_));
 sky130_fd_sc_hd__o31a_1 _20575_ (.A1(_09448_),
    .A2(_09457_),
    .A3(_09903_),
    .B1(_09906_),
    .X(_10339_));
 sky130_fd_sc_hd__a311oi_4 _20576_ (.A1(_10331_),
    .A2(_10332_),
    .A3(net212),
    .B1(_10320_),
    .C1(net326),
    .Y(_10340_));
 sky130_fd_sc_hd__a311o_1 _20577_ (.A1(_10331_),
    .A2(_10332_),
    .A3(net212),
    .B1(_10320_),
    .C1(net326),
    .X(_10341_));
 sky130_fd_sc_hd__a2bb2oi_2 _20578_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_10321_),
    .B2(_10335_),
    .Y(_10342_));
 sky130_fd_sc_hd__o21ai_1 _20579_ (.A1(net361),
    .A2(net345),
    .B1(_10336_),
    .Y(_10343_));
 sky130_fd_sc_hd__o211ai_1 _20580_ (.A1(_09907_),
    .A2(_10337_),
    .B1(_10341_),
    .C1(_10343_),
    .Y(_10345_));
 sky130_fd_sc_hd__o22ai_1 _20581_ (.A1(_09903_),
    .A2(_10338_),
    .B1(_10340_),
    .B2(_10342_),
    .Y(_10346_));
 sky130_fd_sc_hd__nand3_2 _20582_ (.A(_10345_),
    .B(_10346_),
    .C(net211),
    .Y(_10347_));
 sky130_fd_sc_hd__a211o_1 _20583_ (.A1(_10321_),
    .A2(_10335_),
    .B1(_06608_),
    .C1(net237),
    .X(_10348_));
 sky130_fd_sc_hd__o211ai_1 _20584_ (.A1(_09903_),
    .A2(_10338_),
    .B1(_10341_),
    .C1(_10343_),
    .Y(_10349_));
 sky130_fd_sc_hd__o22ai_1 _20585_ (.A1(_09907_),
    .A2(_10337_),
    .B1(_10340_),
    .B2(_10342_),
    .Y(_10350_));
 sky130_fd_sc_hd__nand3_2 _20586_ (.A(_10349_),
    .B(_10350_),
    .C(net211),
    .Y(_10351_));
 sky130_fd_sc_hd__o21ai_4 _20587_ (.A1(net211),
    .A2(_10336_),
    .B1(_10347_),
    .Y(_10352_));
 sky130_fd_sc_hd__o211ai_4 _20588_ (.A1(_10336_),
    .A2(net211),
    .B1(_11309_),
    .C1(_10347_),
    .Y(_10353_));
 sky130_fd_sc_hd__o211ai_4 _20589_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_10348_),
    .C1(_10351_),
    .Y(_10354_));
 sky130_fd_sc_hd__inv_2 _20590_ (.A(_10354_),
    .Y(_10356_));
 sky130_fd_sc_hd__o31a_1 _20591_ (.A1(net365),
    .A2(net362),
    .A3(_09917_),
    .B1(_09584_),
    .X(_10357_));
 sky130_fd_sc_hd__o21ai_1 _20592_ (.A1(_10015_),
    .A2(_09917_),
    .B1(_09925_),
    .Y(_10358_));
 sky130_fd_sc_hd__o2bb2ai_2 _20593_ (.A1_N(_10353_),
    .A2_N(_10354_),
    .B1(_10357_),
    .B2(_09921_),
    .Y(_10359_));
 sky130_fd_sc_hd__o2111ai_4 _20594_ (.A1(_09585_),
    .A2(_09919_),
    .B1(_09922_),
    .C1(_10353_),
    .D1(_10354_),
    .Y(_10360_));
 sky130_fd_sc_hd__a211o_1 _20595_ (.A1(_10348_),
    .A2(_10351_),
    .B1(net230),
    .C1(_06901_),
    .X(_10361_));
 sky130_fd_sc_hd__a31oi_2 _20596_ (.A1(_10353_),
    .A2(_10354_),
    .A3(_10358_),
    .B1(_06904_),
    .Y(_10362_));
 sky130_fd_sc_hd__nand3_4 _20597_ (.A(_10359_),
    .B(_10360_),
    .C(net208),
    .Y(_10363_));
 sky130_fd_sc_hd__o2bb2ai_4 _20598_ (.A1_N(_10362_),
    .A2_N(_10359_),
    .B1(_10352_),
    .B2(net208),
    .Y(_10364_));
 sky130_fd_sc_hd__inv_2 _20599_ (.A(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__a2bb2oi_4 _20600_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_10361_),
    .B2(_10363_),
    .Y(_10367_));
 sky130_fd_sc_hd__o21ai_1 _20601_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_10364_),
    .Y(_10368_));
 sky130_fd_sc_hd__o221a_1 _20602_ (.A1(net365),
    .A2(net362),
    .B1(net208),
    .B2(_10352_),
    .C1(_10363_),
    .X(_10369_));
 sky130_fd_sc_hd__o221ai_4 _20603_ (.A1(net365),
    .A2(net362),
    .B1(net208),
    .B2(_10352_),
    .C1(_10363_),
    .Y(_10370_));
 sky130_fd_sc_hd__a32o_2 _20604_ (.A1(_08874_),
    .A2(_08896_),
    .A3(_09932_),
    .B1(_09935_),
    .B2(_09937_),
    .X(_10371_));
 sky130_fd_sc_hd__o21bai_1 _20605_ (.A1(_10367_),
    .A2(_10369_),
    .B1_N(_10371_),
    .Y(_10372_));
 sky130_fd_sc_hd__o31a_1 _20606_ (.A1(_09927_),
    .A2(_09949_),
    .A3(_10364_),
    .B1(_10371_),
    .X(_10373_));
 sky130_fd_sc_hd__o21ai_2 _20607_ (.A1(_10025_),
    .A2(_10364_),
    .B1(_10371_),
    .Y(_10374_));
 sky130_fd_sc_hd__nand3b_1 _20608_ (.A_N(_10371_),
    .B(_10370_),
    .C(_10368_),
    .Y(_10375_));
 sky130_fd_sc_hd__o21ai_1 _20609_ (.A1(_10367_),
    .A2(_10369_),
    .B1(_10371_),
    .Y(_10376_));
 sky130_fd_sc_hd__o211ai_2 _20610_ (.A1(_07227_),
    .A2(net203),
    .B1(_10375_),
    .C1(_10376_),
    .Y(_10378_));
 sky130_fd_sc_hd__a211o_1 _20611_ (.A1(_10361_),
    .A2(_10363_),
    .B1(_07227_),
    .C1(net203),
    .X(_10379_));
 sky130_fd_sc_hd__o221ai_4 _20612_ (.A1(_07227_),
    .A2(net203),
    .B1(_10367_),
    .B2(_10374_),
    .C1(_10372_),
    .Y(_10380_));
 sky130_fd_sc_hd__o21ai_1 _20613_ (.A1(net185),
    .A2(_10365_),
    .B1(_10380_),
    .Y(_10381_));
 sky130_fd_sc_hd__a211o_2 _20614_ (.A1(_10379_),
    .A2(_10380_),
    .B1(_07544_),
    .C1(net184),
    .X(_10382_));
 sky130_fd_sc_hd__a21oi_2 _20615_ (.A1(_09582_),
    .A2(_09952_),
    .B1(_09953_),
    .Y(_10383_));
 sky130_fd_sc_hd__and3_2 _20616_ (.A(_10380_),
    .B(_08907_),
    .C(_10379_),
    .X(_10384_));
 sky130_fd_sc_hd__o211ai_2 _20617_ (.A1(net185),
    .A2(_10365_),
    .B1(_08907_),
    .C1(_10380_),
    .Y(_10385_));
 sky130_fd_sc_hd__o311a_2 _20618_ (.A1(_07227_),
    .A2(net203),
    .A3(_10364_),
    .B1(_10378_),
    .C1(_08918_),
    .X(_10386_));
 sky130_fd_sc_hd__o211ai_4 _20619_ (.A1(_10364_),
    .A2(net185),
    .B1(_08918_),
    .C1(_10378_),
    .Y(_10387_));
 sky130_fd_sc_hd__o21ai_1 _20620_ (.A1(_09953_),
    .A2(_09955_),
    .B1(_10387_),
    .Y(_10389_));
 sky130_fd_sc_hd__o211a_1 _20621_ (.A1(_09953_),
    .A2(_09955_),
    .B1(_10385_),
    .C1(_10387_),
    .X(_10390_));
 sky130_fd_sc_hd__a21boi_1 _20622_ (.A1(_10385_),
    .A2(_10387_),
    .B1_N(_10383_),
    .Y(_10391_));
 sky130_fd_sc_hd__a21bo_1 _20623_ (.A1(_10385_),
    .A2(_10387_),
    .B1_N(_10383_),
    .X(_10392_));
 sky130_fd_sc_hd__o221ai_4 _20624_ (.A1(_07544_),
    .A2(net184),
    .B1(_10384_),
    .B2(_10389_),
    .C1(_10392_),
    .Y(_10393_));
 sky130_fd_sc_hd__o22ai_2 _20625_ (.A1(_07544_),
    .A2(net184),
    .B1(_10390_),
    .B2(_10391_),
    .Y(_10394_));
 sky130_fd_sc_hd__or3_1 _20626_ (.A(_07544_),
    .B(net184),
    .C(_10381_),
    .X(_10395_));
 sky130_fd_sc_hd__nand2_2 _20627_ (.A(_10382_),
    .B(_10393_),
    .Y(_10396_));
 sky130_fd_sc_hd__a211o_1 _20628_ (.A1(_10382_),
    .A2(_10393_),
    .B1(_07912_),
    .C1(_07914_),
    .X(_10397_));
 sky130_fd_sc_hd__and3_1 _20629_ (.A(_07899_),
    .B(_10394_),
    .C(_10395_),
    .X(_10398_));
 sky130_fd_sc_hd__nand3_4 _20630_ (.A(_07899_),
    .B(_10394_),
    .C(_10395_),
    .Y(_10400_));
 sky130_fd_sc_hd__o311a_1 _20631_ (.A1(_07550_),
    .A2(_10390_),
    .A3(_10391_),
    .B1(_10382_),
    .C1(_07888_),
    .X(_10401_));
 sky130_fd_sc_hd__o211ai_4 _20632_ (.A1(net368),
    .A2(_07866_),
    .B1(_10382_),
    .C1(_10393_),
    .Y(_10402_));
 sky130_fd_sc_hd__o311a_1 _20633_ (.A1(net381),
    .A2(_06310_),
    .A3(_09505_),
    .B1(_09517_),
    .C1(_09968_),
    .X(_10403_));
 sky130_fd_sc_hd__o22a_1 _20634_ (.A1(_09507_),
    .A2(_09516_),
    .B1(_09958_),
    .B2(_09965_),
    .X(_10404_));
 sky130_fd_sc_hd__nor2_1 _20635_ (.A(_09967_),
    .B(_10404_),
    .Y(_10405_));
 sky130_fd_sc_hd__o2bb2ai_2 _20636_ (.A1_N(_10400_),
    .A2_N(_10402_),
    .B1(_10404_),
    .B2(_09967_),
    .Y(_10406_));
 sky130_fd_sc_hd__o2111ai_4 _20637_ (.A1(_09964_),
    .A2(_09966_),
    .B1(_09968_),
    .C1(_10400_),
    .D1(_10402_),
    .Y(_10407_));
 sky130_fd_sc_hd__o2bb2ai_1 _20638_ (.A1_N(_10400_),
    .A2_N(_10402_),
    .B1(_10403_),
    .B2(_09966_),
    .Y(_10408_));
 sky130_fd_sc_hd__o22a_1 _20639_ (.A1(_09967_),
    .A2(_10404_),
    .B1(_10396_),
    .B2(_07899_),
    .X(_10409_));
 sky130_fd_sc_hd__o211ai_1 _20640_ (.A1(_09967_),
    .A2(_10404_),
    .B1(_10402_),
    .C1(_10400_),
    .Y(_10411_));
 sky130_fd_sc_hd__nand3_1 _20641_ (.A(_10408_),
    .B(_10411_),
    .C(net160),
    .Y(_10412_));
 sky130_fd_sc_hd__nand3_1 _20642_ (.A(_10406_),
    .B(_10407_),
    .C(net160),
    .Y(_10413_));
 sky130_fd_sc_hd__o311a_2 _20643_ (.A1(_07550_),
    .A2(_10390_),
    .A3(_10391_),
    .B1(_07917_),
    .C1(_10382_),
    .X(_10414_));
 sky130_fd_sc_hd__a31o_1 _20644_ (.A1(_10406_),
    .A2(_10407_),
    .A3(net160),
    .B1(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__a31oi_4 _20645_ (.A1(_10406_),
    .A2(_10407_),
    .A3(net160),
    .B1(_10414_),
    .Y(_10416_));
 sky130_fd_sc_hd__and3_1 _20646_ (.A(_10412_),
    .B(_07033_),
    .C(_10397_),
    .X(_10417_));
 sky130_fd_sc_hd__o211ai_2 _20647_ (.A1(_06989_),
    .A2(net375),
    .B1(_10397_),
    .C1(_10412_),
    .Y(_10418_));
 sky130_fd_sc_hd__o211a_1 _20648_ (.A1(_10396_),
    .A2(net160),
    .B1(_07044_),
    .C1(_10413_),
    .X(_10419_));
 sky130_fd_sc_hd__o2111ai_4 _20649_ (.A1(_10396_),
    .A2(net160),
    .B1(_07022_),
    .C1(net376),
    .D1(_10413_),
    .Y(_10420_));
 sky130_fd_sc_hd__o211a_1 _20650_ (.A1(_09974_),
    .A2(_09981_),
    .B1(_10418_),
    .C1(_10420_),
    .X(_10422_));
 sky130_fd_sc_hd__a21oi_2 _20651_ (.A1(_10418_),
    .A2(_10420_),
    .B1(_10019_),
    .Y(_10423_));
 sky130_fd_sc_hd__a21o_1 _20652_ (.A1(_10418_),
    .A2(_10420_),
    .B1(_10019_),
    .X(_10424_));
 sky130_fd_sc_hd__o22ai_2 _20653_ (.A1(net180),
    .A2(_08298_),
    .B1(_10422_),
    .B2(_10423_),
    .Y(_10425_));
 sky130_fd_sc_hd__a311o_1 _20654_ (.A1(_10406_),
    .A2(_10407_),
    .A3(net160),
    .B1(_10414_),
    .C1(_08300_),
    .X(_10426_));
 sky130_fd_sc_hd__nand3b_1 _20655_ (.A_N(_10422_),
    .B(_10424_),
    .C(_08300_),
    .Y(_10427_));
 sky130_fd_sc_hd__o31a_1 _20656_ (.A1(_08301_),
    .A2(_10422_),
    .A3(_10423_),
    .B1(_10426_),
    .X(_10428_));
 sky130_fd_sc_hd__or3_2 _20657_ (.A(net158),
    .B(_08712_),
    .C(_10428_),
    .X(_10429_));
 sky130_fd_sc_hd__o2111ai_4 _20658_ (.A1(_10416_),
    .A2(_08300_),
    .B1(_06321_),
    .C1(_06300_),
    .D1(_10425_),
    .Y(_10430_));
 sky130_fd_sc_hd__o311a_1 _20659_ (.A1(_08301_),
    .A2(_10422_),
    .A3(_10423_),
    .B1(_10426_),
    .C1(_06332_),
    .X(_10431_));
 sky130_fd_sc_hd__o221ai_2 _20660_ (.A1(net381),
    .A2(_06310_),
    .B1(_08300_),
    .B2(_10415_),
    .C1(_10427_),
    .Y(_10433_));
 sky130_fd_sc_hd__a21oi_1 _20661_ (.A1(_05862_),
    .A2(_09988_),
    .B1(_09990_),
    .Y(_10434_));
 sky130_fd_sc_hd__a32oi_4 _20662_ (.A1(net406),
    .A2(_05840_),
    .A3(_09990_),
    .B1(_09991_),
    .B2(_09988_),
    .Y(_10435_));
 sky130_fd_sc_hd__o2bb2ai_2 _20663_ (.A1_N(_10430_),
    .A2_N(_10433_),
    .B1(_10434_),
    .B2(_09996_),
    .Y(_10436_));
 sky130_fd_sc_hd__a31oi_1 _20664_ (.A1(_10427_),
    .A2(_06332_),
    .A3(_10426_),
    .B1(_10435_),
    .Y(_10437_));
 sky130_fd_sc_hd__o21ai_2 _20665_ (.A1(_06332_),
    .A2(_10428_),
    .B1(_10437_),
    .Y(_10438_));
 sky130_fd_sc_hd__o211ai_4 _20666_ (.A1(net158),
    .A2(_08712_),
    .B1(_10436_),
    .C1(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__a22oi_2 _20667_ (.A1(_08710_),
    .A2(_08713_),
    .B1(_10436_),
    .B2(_10438_),
    .Y(_10440_));
 sky130_fd_sc_hd__o311a_1 _20668_ (.A1(_08301_),
    .A2(_10422_),
    .A3(_10423_),
    .B1(_10426_),
    .C1(_08715_),
    .X(_10441_));
 sky130_fd_sc_hd__o311ai_4 _20669_ (.A1(_09994_),
    .A2(_09987_),
    .A3(_09985_),
    .B1(_09999_),
    .C1(_09995_),
    .Y(_10442_));
 sky130_fd_sc_hd__o31ai_2 _20670_ (.A1(_05545_),
    .A2(_09540_),
    .A3(_09543_),
    .B1(_10442_),
    .Y(_10444_));
 sky130_fd_sc_hd__and3_2 _20671_ (.A(_10442_),
    .B(_05851_),
    .C(_10000_),
    .X(_10445_));
 sky130_fd_sc_hd__a22o_2 _20672_ (.A1(net395),
    .A2(_05796_),
    .B1(_10000_),
    .B2(_10442_),
    .X(_10446_));
 sky130_fd_sc_hd__a2bb2o_1 _20673_ (.A1_N(_09120_),
    .A2_N(_09121_),
    .B1(_10444_),
    .B2(_05862_),
    .X(_10447_));
 sky130_fd_sc_hd__o311ai_4 _20674_ (.A1(_05763_),
    .A2(_05785_),
    .A3(_10444_),
    .B1(_10446_),
    .C1(_09125_),
    .Y(_10448_));
 sky130_fd_sc_hd__o221a_1 _20675_ (.A1(_08714_),
    .A2(_10428_),
    .B1(_10445_),
    .B2(_10447_),
    .C1(_10439_),
    .X(_10449_));
 sky130_fd_sc_hd__o221ai_2 _20676_ (.A1(_08714_),
    .A2(_10428_),
    .B1(_10445_),
    .B2(_10447_),
    .C1(_10439_),
    .Y(_10450_));
 sky130_fd_sc_hd__a21oi_1 _20677_ (.A1(_10429_),
    .A2(_10439_),
    .B1(_10448_),
    .Y(_10451_));
 sky130_fd_sc_hd__o31a_1 _20678_ (.A1(_10448_),
    .A2(_10441_),
    .A3(_10440_),
    .B1(_10450_),
    .X(_10452_));
 sky130_fd_sc_hd__o21ai_1 _20679_ (.A1(_09549_),
    .A2(_10006_),
    .B1(_10008_),
    .Y(_10453_));
 sky130_fd_sc_hd__o221ai_4 _20680_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_09549_),
    .B2(_10006_),
    .C1(_10008_),
    .Y(_10455_));
 sky130_fd_sc_hd__o21ai_1 _20681_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_10453_),
    .Y(_10456_));
 sky130_fd_sc_hd__a21oi_1 _20682_ (.A1(_05556_),
    .A2(_10453_),
    .B1(_09562_),
    .Y(_10457_));
 sky130_fd_sc_hd__o211ai_1 _20683_ (.A1(_09553_),
    .A2(net155),
    .B1(_10455_),
    .C1(_10456_),
    .Y(_10458_));
 sky130_fd_sc_hd__nand3_2 _20684_ (.A(_10452_),
    .B(_10455_),
    .C(_10457_),
    .Y(_10459_));
 sky130_fd_sc_hd__o21ai_2 _20685_ (.A1(_10449_),
    .A2(_10451_),
    .B1(_10458_),
    .Y(_10460_));
 sky130_fd_sc_hd__nand2_1 _20686_ (.A(_10459_),
    .B(_10460_),
    .Y(_10461_));
 sky130_fd_sc_hd__a21oi_2 _20687_ (.A1(_10459_),
    .A2(_10460_),
    .B1(_05239_),
    .Y(_10462_));
 sky130_fd_sc_hd__nand4_2 _20688_ (.A(_05207_),
    .B(_05229_),
    .C(_10459_),
    .D(_10460_),
    .Y(_10463_));
 sky130_fd_sc_hd__a41o_1 _20689_ (.A1(_05207_),
    .A2(_05229_),
    .A3(_10459_),
    .A4(_10460_),
    .B1(_10462_),
    .X(_10464_));
 sky130_fd_sc_hd__and4b_1 _20690_ (.A_N(_10462_),
    .B(_10463_),
    .C(net1),
    .D(_10012_),
    .X(_10466_));
 sky130_fd_sc_hd__a22o_1 _20691_ (.A1(_09572_),
    .A2(_09574_),
    .B1(_10013_),
    .B2(_10464_),
    .X(_10467_));
 sky130_fd_sc_hd__o22ai_1 _20692_ (.A1(_09579_),
    .A2(_10461_),
    .B1(_10466_),
    .B2(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__o32a_1 _20693_ (.A1(_09571_),
    .A2(_09573_),
    .A3(_10461_),
    .B1(_10466_),
    .B2(_10467_),
    .X(_10469_));
 sky130_fd_sc_hd__nor2_1 _20694_ (.A(_03289_),
    .B(_10469_),
    .Y(_10470_));
 sky130_fd_sc_hd__nand2_1 _20695_ (.A(net1),
    .B(_10468_),
    .Y(_10471_));
 sky130_fd_sc_hd__o221a_1 _20696_ (.A1(_09579_),
    .A2(_10461_),
    .B1(_10466_),
    .B2(_10467_),
    .C1(_03289_),
    .X(_10472_));
 sky130_fd_sc_hd__or4_4 _20697_ (.A(net50),
    .B(net51),
    .C(net52),
    .D(_09118_),
    .X(_10473_));
 sky130_fd_sc_hd__and3b_4 _20698_ (.A_N(net53),
    .B(_10473_),
    .C(net409),
    .X(_10474_));
 sky130_fd_sc_hd__a21boi_4 _20699_ (.A1(_10473_),
    .A2(net409),
    .B1_N(net53),
    .Y(_10475_));
 sky130_fd_sc_hd__a21oi_4 _20700_ (.A1(_10473_),
    .A2(net409),
    .B1(net53),
    .Y(_10477_));
 sky130_fd_sc_hd__o311a_4 _20701_ (.A1(net51),
    .A2(net52),
    .A3(_09552_),
    .B1(net53),
    .C1(net409),
    .X(_10478_));
 sky130_fd_sc_hd__nor2_8 _20702_ (.A(_10474_),
    .B(net138),
    .Y(_10479_));
 sky130_fd_sc_hd__nor2_8 _20703_ (.A(_10477_),
    .B(_10478_),
    .Y(_10480_));
 sky130_fd_sc_hd__or3_1 _20704_ (.A(_10474_),
    .B(net138),
    .C(_10469_),
    .X(_10481_));
 sky130_fd_sc_hd__o31a_1 _20705_ (.A1(_10470_),
    .A2(_10472_),
    .A3(_10479_),
    .B1(_10481_),
    .X(_10482_));
 sky130_fd_sc_hd__xor2_1 _20706_ (.A(_10018_),
    .B(_10482_),
    .X(net85));
 sky130_fd_sc_hd__and4_1 _20707_ (.A(_09130_),
    .B(_09565_),
    .C(_10017_),
    .D(_10482_),
    .X(_10483_));
 sky130_fd_sc_hd__o21ai_2 _20708_ (.A1(_10431_),
    .A2(_10435_),
    .B1(_10430_),
    .Y(_10484_));
 sky130_fd_sc_hd__or4_4 _20709_ (.A(net19),
    .B(net20),
    .C(net21),
    .D(_09133_),
    .X(_10485_));
 sky130_fd_sc_hd__and3b_4 _20710_ (.A_N(net22),
    .B(_10485_),
    .C(net410),
    .X(_10487_));
 sky130_fd_sc_hd__a21boi_4 _20711_ (.A1(_10485_),
    .A2(net410),
    .B1_N(net22),
    .Y(_10488_));
 sky130_fd_sc_hd__a21oi_4 _20712_ (.A1(_10485_),
    .A2(net410),
    .B1(net22),
    .Y(_10489_));
 sky130_fd_sc_hd__o311a_4 _20713_ (.A1(net20),
    .A2(net21),
    .A3(_09586_),
    .B1(net22),
    .C1(net410),
    .X(_10490_));
 sky130_fd_sc_hd__nor2_8 _20714_ (.A(_10487_),
    .B(net165),
    .Y(_10491_));
 sky130_fd_sc_hd__nor2_8 _20715_ (.A(net164),
    .B(_10490_),
    .Y(_10492_));
 sky130_fd_sc_hd__o221a_2 _20716_ (.A1(_05130_),
    .A2(_05152_),
    .B1(_10487_),
    .B2(net166),
    .C1(net33),
    .X(_10493_));
 sky130_fd_sc_hd__nor4_1 _20717_ (.A(_08745_),
    .B(_09145_),
    .C(_09599_),
    .D(_10032_),
    .Y(_10494_));
 sky130_fd_sc_hd__or4_1 _20718_ (.A(_08745_),
    .B(_09145_),
    .C(_09599_),
    .D(_10032_),
    .X(_10495_));
 sky130_fd_sc_hd__nand2_1 _20719_ (.A(_08740_),
    .B(_10494_),
    .Y(_10496_));
 sky130_fd_sc_hd__a31o_1 _20720_ (.A1(net33),
    .A2(_09595_),
    .A3(net151),
    .B1(_10494_),
    .X(_10498_));
 sky130_fd_sc_hd__o21bai_4 _20721_ (.A1(_10032_),
    .A2(_10034_),
    .B1_N(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__and3_1 _20722_ (.A(_10492_),
    .B(net33),
    .C(net151),
    .X(_10500_));
 sky130_fd_sc_hd__or4_1 _20723_ (.A(_10489_),
    .B(_03178_),
    .C(net153),
    .D(_10490_),
    .X(_10501_));
 sky130_fd_sc_hd__o32a_1 _20724_ (.A1(_03178_),
    .A2(_10489_),
    .A3(_10490_),
    .B1(_10023_),
    .B2(_10024_),
    .X(_10502_));
 sky130_fd_sc_hd__a21oi_1 _20725_ (.A1(_10028_),
    .A2(_10492_),
    .B1(_10502_),
    .Y(_10503_));
 sky130_fd_sc_hd__o2bb2ai_4 _20726_ (.A1_N(_10496_),
    .A2_N(_10499_),
    .B1(_10500_),
    .B2(_10502_),
    .Y(_10504_));
 sky130_fd_sc_hd__o211ai_4 _20727_ (.A1(_08739_),
    .A2(_10495_),
    .B1(_10503_),
    .C1(_10499_),
    .Y(_10505_));
 sky130_fd_sc_hd__nand2_1 _20728_ (.A(_10504_),
    .B(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__a22o_1 _20729_ (.A1(_05141_),
    .A2(_05163_),
    .B1(_10492_),
    .B2(net33),
    .X(_10507_));
 sky130_fd_sc_hd__a31oi_4 _20730_ (.A1(_10504_),
    .A2(_10505_),
    .A3(net405),
    .B1(_10493_),
    .Y(_10509_));
 sky130_fd_sc_hd__a31o_1 _20731_ (.A1(_10504_),
    .A2(_10505_),
    .A3(net405),
    .B1(_10493_),
    .X(_10510_));
 sky130_fd_sc_hd__or3_1 _20732_ (.A(_05348_),
    .B(net401),
    .C(_10509_),
    .X(_10511_));
 sky130_fd_sc_hd__a311oi_4 _20733_ (.A1(_10504_),
    .A2(_10505_),
    .A3(net405),
    .B1(_09595_),
    .C1(_10493_),
    .Y(_10512_));
 sky130_fd_sc_hd__a311o_1 _20734_ (.A1(_10504_),
    .A2(_10505_),
    .A3(net405),
    .B1(_09595_),
    .C1(_10493_),
    .X(_10513_));
 sky130_fd_sc_hd__a22oi_1 _20735_ (.A1(_09589_),
    .A2(_09591_),
    .B1(_10506_),
    .B2(net405),
    .Y(_10514_));
 sky130_fd_sc_hd__a21oi_1 _20736_ (.A1(_09589_),
    .A2(_09591_),
    .B1(_10509_),
    .Y(_10515_));
 sky130_fd_sc_hd__o21ai_2 _20737_ (.A1(_09588_),
    .A2(net187),
    .B1(_10510_),
    .Y(_10516_));
 sky130_fd_sc_hd__a21oi_1 _20738_ (.A1(_10514_),
    .A2(_10507_),
    .B1(_10512_),
    .Y(_10517_));
 sky130_fd_sc_hd__o221ai_4 _20739_ (.A1(net177),
    .A2(_09606_),
    .B1(_09612_),
    .B2(_09616_),
    .C1(_10044_),
    .Y(_10518_));
 sky130_fd_sc_hd__o2111ai_4 _20740_ (.A1(net173),
    .A2(_10041_),
    .B1(_10513_),
    .C1(_10516_),
    .D1(_10518_),
    .Y(_10520_));
 sky130_fd_sc_hd__o21ai_1 _20741_ (.A1(_10512_),
    .A2(_10515_),
    .B1(_10044_),
    .Y(_10521_));
 sky130_fd_sc_hd__o211ai_4 _20742_ (.A1(_10049_),
    .A2(_10521_),
    .B1(_10520_),
    .C1(_05403_),
    .Y(_10522_));
 sky130_fd_sc_hd__o21a_2 _20743_ (.A1(_05403_),
    .A2(_10509_),
    .B1(_10522_),
    .X(_10523_));
 sky130_fd_sc_hd__o21ai_2 _20744_ (.A1(_05403_),
    .A2(_10509_),
    .B1(_10522_),
    .Y(_10524_));
 sky130_fd_sc_hd__and3_1 _20745_ (.A(_05731_),
    .B(_10511_),
    .C(_10522_),
    .X(_10525_));
 sky130_fd_sc_hd__o32ai_1 _20746_ (.A1(_08728_),
    .A2(net195),
    .A3(_10054_),
    .B1(_10064_),
    .B2(_10065_),
    .Y(_10526_));
 sky130_fd_sc_hd__a2bb2o_1 _20747_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_10511_),
    .B2(_10522_),
    .X(_10527_));
 sky130_fd_sc_hd__o211ai_4 _20748_ (.A1(_05403_),
    .A2(_10509_),
    .B1(net174),
    .C1(_10522_),
    .Y(_10528_));
 sky130_fd_sc_hd__nand2_1 _20749_ (.A(_10527_),
    .B(_10528_),
    .Y(_10529_));
 sky130_fd_sc_hd__a21oi_2 _20750_ (.A1(_10060_),
    .A2(_10067_),
    .B1(_10529_),
    .Y(_10531_));
 sky130_fd_sc_hd__nand3_1 _20751_ (.A(_10526_),
    .B(_10527_),
    .C(_10528_),
    .Y(_10532_));
 sky130_fd_sc_hd__o311a_1 _20752_ (.A1(_08728_),
    .A2(net195),
    .A3(_10054_),
    .B1(_10067_),
    .C1(_10529_),
    .X(_10533_));
 sky130_fd_sc_hd__o211ai_1 _20753_ (.A1(_10064_),
    .A2(_10065_),
    .B1(_10529_),
    .C1(_10060_),
    .Y(_10534_));
 sky130_fd_sc_hd__o22a_1 _20754_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_10531_),
    .B2(_10533_),
    .X(_10535_));
 sky130_fd_sc_hd__o22ai_2 _20755_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_10531_),
    .B2(_10533_),
    .Y(_10536_));
 sky130_fd_sc_hd__or3_1 _20756_ (.A(_05676_),
    .B(_05698_),
    .C(_10523_),
    .X(_10537_));
 sky130_fd_sc_hd__nand3_1 _20757_ (.A(_10532_),
    .B(_10534_),
    .C(net358),
    .Y(_10538_));
 sky130_fd_sc_hd__a31o_2 _20758_ (.A1(_05731_),
    .A2(_10511_),
    .A3(_10522_),
    .B1(_10535_),
    .X(_10539_));
 sky130_fd_sc_hd__or4_4 _20759_ (.A(_06793_),
    .B(_06815_),
    .C(_10525_),
    .D(_10535_),
    .X(_10540_));
 sky130_fd_sc_hd__a2bb2oi_1 _20760_ (.A1_N(_08724_),
    .A2_N(_08726_),
    .B1(_10537_),
    .B2(_10538_),
    .Y(_10542_));
 sky130_fd_sc_hd__o211ai_4 _20761_ (.A1(_10524_),
    .A2(net358),
    .B1(net175),
    .C1(_10536_),
    .Y(_10543_));
 sky130_fd_sc_hd__a31oi_1 _20762_ (.A1(_10532_),
    .A2(_10534_),
    .A3(net358),
    .B1(net175),
    .Y(_10544_));
 sky130_fd_sc_hd__o211ai_2 _20763_ (.A1(net358),
    .A2(_10523_),
    .B1(net177),
    .C1(_10538_),
    .Y(_10545_));
 sky130_fd_sc_hd__a21oi_2 _20764_ (.A1(_10537_),
    .A2(_10544_),
    .B1(_10542_),
    .Y(_10546_));
 sky130_fd_sc_hd__nand2_4 _20765_ (.A(_10543_),
    .B(_10545_),
    .Y(_10547_));
 sky130_fd_sc_hd__a31oi_4 _20766_ (.A1(_10088_),
    .A2(_10090_),
    .A3(_10081_),
    .B1(_10075_),
    .Y(_10548_));
 sky130_fd_sc_hd__o22ai_2 _20767_ (.A1(net199),
    .A2(_10072_),
    .B1(_10094_),
    .B2(_10087_),
    .Y(_10549_));
 sky130_fd_sc_hd__a21oi_1 _20768_ (.A1(_10076_),
    .A2(_10095_),
    .B1(_10547_),
    .Y(_10550_));
 sky130_fd_sc_hd__nand2_1 _20769_ (.A(_10549_),
    .B(_10546_),
    .Y(_10551_));
 sky130_fd_sc_hd__o211ai_2 _20770_ (.A1(net199),
    .A2(_10072_),
    .B1(_10095_),
    .C1(_10547_),
    .Y(_10553_));
 sky130_fd_sc_hd__o22ai_2 _20771_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_10546_),
    .B2(_10549_),
    .Y(_10554_));
 sky130_fd_sc_hd__nand3_2 _20772_ (.A(_10551_),
    .B(_10553_),
    .C(net357),
    .Y(_10555_));
 sky130_fd_sc_hd__o22a_2 _20773_ (.A1(net357),
    .A2(_10539_),
    .B1(_10550_),
    .B2(_10554_),
    .X(_10556_));
 sky130_fd_sc_hd__o22ai_2 _20774_ (.A1(net357),
    .A2(_10539_),
    .B1(_10550_),
    .B2(_10554_),
    .Y(_10557_));
 sky130_fd_sc_hd__a21oi_2 _20775_ (.A1(_10540_),
    .A2(_10555_),
    .B1(net355),
    .Y(_10558_));
 sky130_fd_sc_hd__inv_2 _20776_ (.A(_10558_),
    .Y(_10559_));
 sky130_fd_sc_hd__a2bb2oi_4 _20777_ (.A1_N(_08307_),
    .A2_N(_08309_),
    .B1(_10540_),
    .B2(_10555_),
    .Y(_10560_));
 sky130_fd_sc_hd__o21ai_1 _20778_ (.A1(_08307_),
    .A2(_08309_),
    .B1(_10557_),
    .Y(_10561_));
 sky130_fd_sc_hd__a31oi_2 _20779_ (.A1(_10551_),
    .A2(_10553_),
    .A3(net357),
    .B1(net198),
    .Y(_10562_));
 sky130_fd_sc_hd__o221a_1 _20780_ (.A1(net357),
    .A2(_10539_),
    .B1(_10550_),
    .B2(_10554_),
    .C1(net199),
    .X(_10564_));
 sky130_fd_sc_hd__o221ai_1 _20781_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_10539_),
    .B2(net357),
    .C1(_10555_),
    .Y(_10565_));
 sky130_fd_sc_hd__a21oi_4 _20782_ (.A1(_10540_),
    .A2(_10562_),
    .B1(_10560_),
    .Y(_10566_));
 sky130_fd_sc_hd__nand2_1 _20783_ (.A(_10561_),
    .B(_10565_),
    .Y(_10567_));
 sky130_fd_sc_hd__o211a_1 _20784_ (.A1(_09205_),
    .A2(_09215_),
    .B1(_08805_),
    .C1(_09213_),
    .X(_10568_));
 sky130_fd_sc_hd__nand3_1 _20785_ (.A(_10568_),
    .B(_09677_),
    .C(_09673_),
    .Y(_10569_));
 sky130_fd_sc_hd__o211ai_4 _20786_ (.A1(_09679_),
    .A2(_09680_),
    .B1(_10569_),
    .C1(_09673_),
    .Y(_10570_));
 sky130_fd_sc_hd__a32oi_4 _20787_ (.A1(_09678_),
    .A2(_10568_),
    .A3(_08814_),
    .B1(_10101_),
    .B2(_07935_),
    .Y(_10571_));
 sky130_fd_sc_hd__nand2_1 _20788_ (.A(_10571_),
    .B(_10570_),
    .Y(_10572_));
 sky130_fd_sc_hd__a2bb2oi_4 _20789_ (.A1_N(_07935_),
    .A2_N(_10101_),
    .B1(_10570_),
    .B2(_10571_),
    .Y(_10573_));
 sky130_fd_sc_hd__o2bb2ai_2 _20790_ (.A1_N(_10570_),
    .A2_N(_10571_),
    .B1(_07935_),
    .B2(_10101_),
    .Y(_10575_));
 sky130_fd_sc_hd__o221a_2 _20791_ (.A1(_07935_),
    .A2(_10101_),
    .B1(_10560_),
    .B2(_10564_),
    .C1(_10572_),
    .X(_10576_));
 sky130_fd_sc_hd__o221ai_4 _20792_ (.A1(_07935_),
    .A2(_10101_),
    .B1(_10560_),
    .B2(_10564_),
    .C1(_10572_),
    .Y(_10577_));
 sky130_fd_sc_hd__nand2_2 _20793_ (.A(_10575_),
    .B(_10566_),
    .Y(_10578_));
 sky130_fd_sc_hd__o22ai_4 _20794_ (.A1(_07691_),
    .A2(net371),
    .B1(_10567_),
    .B2(_10573_),
    .Y(_10579_));
 sky130_fd_sc_hd__nand3_1 _20795_ (.A(_10578_),
    .B(net355),
    .C(_10577_),
    .Y(_10580_));
 sky130_fd_sc_hd__o22a_2 _20796_ (.A1(net355),
    .A2(_10556_),
    .B1(_10576_),
    .B2(_10579_),
    .X(_10581_));
 sky130_fd_sc_hd__o22ai_2 _20797_ (.A1(net355),
    .A2(_10556_),
    .B1(_10576_),
    .B2(_10579_),
    .Y(_10582_));
 sky130_fd_sc_hd__or3_2 _20798_ (.A(_08678_),
    .B(_08700_),
    .C(_10581_),
    .X(_10583_));
 sky130_fd_sc_hd__a21oi_1 _20799_ (.A1(_09692_),
    .A2(_10127_),
    .B1(_10120_),
    .Y(_10584_));
 sky130_fd_sc_hd__o211ai_1 _20800_ (.A1(net222),
    .A2(_09688_),
    .B1(_10125_),
    .C1(_10127_),
    .Y(_10586_));
 sky130_fd_sc_hd__o21ai_1 _20801_ (.A1(_07564_),
    .A2(_10119_),
    .B1(_10586_),
    .Y(_10587_));
 sky130_fd_sc_hd__a31oi_4 _20802_ (.A1(_09692_),
    .A2(_10125_),
    .A3(_10127_),
    .B1(_10120_),
    .Y(_10588_));
 sky130_fd_sc_hd__a311oi_4 _20803_ (.A1(_10578_),
    .A2(net355),
    .A3(_10577_),
    .B1(_07936_),
    .C1(_10558_),
    .Y(_10589_));
 sky130_fd_sc_hd__o221ai_4 _20804_ (.A1(net355),
    .A2(_10556_),
    .B1(_10576_),
    .B2(_10579_),
    .C1(_07935_),
    .Y(_10590_));
 sky130_fd_sc_hd__a2bb2oi_2 _20805_ (.A1_N(_07928_),
    .A2_N(_07930_),
    .B1(_10559_),
    .B2(_10580_),
    .Y(_10591_));
 sky130_fd_sc_hd__o21ai_4 _20806_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_10582_),
    .Y(_10592_));
 sky130_fd_sc_hd__nor2_1 _20807_ (.A(_10589_),
    .B(_10591_),
    .Y(_10593_));
 sky130_fd_sc_hd__nand3_2 _20808_ (.A(_10592_),
    .B(_10587_),
    .C(_10590_),
    .Y(_10594_));
 sky130_fd_sc_hd__o22ai_2 _20809_ (.A1(_10123_),
    .A2(_10584_),
    .B1(_10589_),
    .B2(_10591_),
    .Y(_10595_));
 sky130_fd_sc_hd__o211ai_4 _20810_ (.A1(_08678_),
    .A2(_08700_),
    .B1(_10594_),
    .C1(_10595_),
    .Y(_10597_));
 sky130_fd_sc_hd__o21ai_4 _20811_ (.A1(net338),
    .A2(_10581_),
    .B1(_10597_),
    .Y(_10598_));
 sky130_fd_sc_hd__a2bb2oi_4 _20812_ (.A1_N(_07555_),
    .A2_N(net218),
    .B1(_10583_),
    .B2(_10597_),
    .Y(_10599_));
 sky130_fd_sc_hd__a22o_1 _20813_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_10583_),
    .B2(_10597_),
    .X(_10600_));
 sky130_fd_sc_hd__o211a_2 _20814_ (.A1(net338),
    .A2(_10581_),
    .B1(_07564_),
    .C1(_10597_),
    .X(_10601_));
 sky130_fd_sc_hd__o211ai_4 _20815_ (.A1(net338),
    .A2(_10581_),
    .B1(_07564_),
    .C1(_10597_),
    .Y(_10602_));
 sky130_fd_sc_hd__o211a_1 _20816_ (.A1(_10136_),
    .A2(net224),
    .B1(_09709_),
    .C1(_10142_),
    .X(_10603_));
 sky130_fd_sc_hd__o211ai_4 _20817_ (.A1(_10136_),
    .A2(net224),
    .B1(_09709_),
    .C1(_10142_),
    .Y(_10604_));
 sky130_fd_sc_hd__nand4_2 _20818_ (.A(_10138_),
    .B(_10144_),
    .C(_10600_),
    .D(_10602_),
    .Y(_10605_));
 sky130_fd_sc_hd__o221ai_4 _20819_ (.A1(net222),
    .A2(_10134_),
    .B1(_10599_),
    .B2(_10601_),
    .C1(_10604_),
    .Y(_10606_));
 sky130_fd_sc_hd__o211ai_4 _20820_ (.A1(net351),
    .A2(_09807_),
    .B1(_10605_),
    .C1(_10606_),
    .Y(_10608_));
 sky130_fd_sc_hd__a211o_1 _20821_ (.A1(_10583_),
    .A2(_10597_),
    .B1(net351),
    .C1(_09807_),
    .X(_10609_));
 sky130_fd_sc_hd__o22ai_1 _20822_ (.A1(_10599_),
    .A2(_10601_),
    .B1(_10603_),
    .B2(_10139_),
    .Y(_10610_));
 sky130_fd_sc_hd__o2111ai_1 _20823_ (.A1(_10134_),
    .A2(net222),
    .B1(_10602_),
    .C1(_10600_),
    .D1(_10604_),
    .Y(_10611_));
 sky130_fd_sc_hd__o211ai_2 _20824_ (.A1(net351),
    .A2(_09807_),
    .B1(_10610_),
    .C1(_10611_),
    .Y(_10612_));
 sky130_fd_sc_hd__o21a_2 _20825_ (.A1(net335),
    .A2(_10598_),
    .B1(_10608_),
    .X(_10613_));
 sky130_fd_sc_hd__o21ai_4 _20826_ (.A1(net335),
    .A2(_10598_),
    .B1(_10608_),
    .Y(_10614_));
 sky130_fd_sc_hd__o211ai_4 _20827_ (.A1(_10598_),
    .A2(net335),
    .B1(net222),
    .C1(_10608_),
    .Y(_10615_));
 sky130_fd_sc_hd__o211ai_4 _20828_ (.A1(_07244_),
    .A2(_07245_),
    .B1(_10609_),
    .C1(_10612_),
    .Y(_10616_));
 sky130_fd_sc_hd__nand2_1 _20829_ (.A(_10615_),
    .B(_10616_),
    .Y(_10617_));
 sky130_fd_sc_hd__o21ai_1 _20830_ (.A1(net225),
    .A2(_10148_),
    .B1(_10162_),
    .Y(_10619_));
 sky130_fd_sc_hd__o221ai_4 _20831_ (.A1(net225),
    .A2(_10148_),
    .B1(_08455_),
    .B2(_10161_),
    .C1(_10164_),
    .Y(_10620_));
 sky130_fd_sc_hd__o22ai_1 _20832_ (.A1(net227),
    .A2(_10149_),
    .B1(_10619_),
    .B2(_10163_),
    .Y(_10621_));
 sky130_fd_sc_hd__o211ai_2 _20833_ (.A1(net227),
    .A2(_10149_),
    .B1(_10173_),
    .C1(_10617_),
    .Y(_10622_));
 sky130_fd_sc_hd__nand3_2 _20834_ (.A(_10621_),
    .B(_10616_),
    .C(_10615_),
    .Y(_10623_));
 sky130_fd_sc_hd__o211ai_4 _20835_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_10622_),
    .C1(_10623_),
    .Y(_10624_));
 sky130_fd_sc_hd__or3_2 _20836_ (.A(_11046_),
    .B(_11057_),
    .C(_10614_),
    .X(_10625_));
 sky130_fd_sc_hd__o31a_4 _20837_ (.A1(_11046_),
    .A2(_11057_),
    .A3(_10614_),
    .B1(_10624_),
    .X(_10626_));
 sky130_fd_sc_hd__a21oi_2 _20838_ (.A1(_10624_),
    .A2(_10625_),
    .B1(net311),
    .Y(_10627_));
 sky130_fd_sc_hd__or3_1 _20839_ (.A(_12670_),
    .B(net327),
    .C(_10626_),
    .X(_10628_));
 sky130_fd_sc_hd__a22oi_4 _20840_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_10624_),
    .B2(_10625_),
    .Y(_10630_));
 sky130_fd_sc_hd__a22o_1 _20841_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_10624_),
    .B2(_10625_),
    .X(_10631_));
 sky130_fd_sc_hd__a31oi_1 _20842_ (.A1(_10622_),
    .A2(_10623_),
    .A3(net332),
    .B1(net225),
    .Y(_10632_));
 sky130_fd_sc_hd__o221ai_4 _20843_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_10614_),
    .B2(net333),
    .C1(_10624_),
    .Y(_10633_));
 sky130_fd_sc_hd__a21oi_2 _20844_ (.A1(_10625_),
    .A2(_10632_),
    .B1(_10630_),
    .Y(_10634_));
 sky130_fd_sc_hd__nand3_1 _20845_ (.A(_09288_),
    .B(_09290_),
    .C(_08875_),
    .Y(_10635_));
 sky130_fd_sc_hd__a211oi_4 _20846_ (.A1(_09729_),
    .A2(_09743_),
    .B1(_10635_),
    .C1(_09747_),
    .Y(_10636_));
 sky130_fd_sc_hd__nand2_1 _20847_ (.A(_10180_),
    .B(_10636_),
    .Y(_10637_));
 sky130_fd_sc_hd__a21oi_1 _20848_ (.A1(_10180_),
    .A2(_10636_),
    .B1(_10181_),
    .Y(_10638_));
 sky130_fd_sc_hd__o211ai_4 _20849_ (.A1(_10185_),
    .A2(_10178_),
    .B1(_10182_),
    .C1(_10637_),
    .Y(_10639_));
 sky130_fd_sc_hd__nand3_2 _20850_ (.A(_10180_),
    .B(_10182_),
    .C(_10636_),
    .Y(_10641_));
 sky130_fd_sc_hd__o211ai_2 _20851_ (.A1(_08881_),
    .A2(_08884_),
    .B1(_10636_),
    .C1(_10182_),
    .Y(_10642_));
 sky130_fd_sc_hd__nand4b_1 _20852_ (.A_N(_08886_),
    .B(_10180_),
    .C(_10182_),
    .D(_10636_),
    .Y(_10643_));
 sky130_fd_sc_hd__a2bb2oi_4 _20853_ (.A1_N(_10178_),
    .A2_N(_10642_),
    .B1(_10187_),
    .B2(_10638_),
    .Y(_10644_));
 sky130_fd_sc_hd__o2111a_2 _20854_ (.A1(_10641_),
    .A2(_08886_),
    .B1(_10633_),
    .C1(_10639_),
    .D1(_10631_),
    .X(_10645_));
 sky130_fd_sc_hd__o2111ai_4 _20855_ (.A1(_10641_),
    .A2(_08886_),
    .B1(_10633_),
    .C1(_10639_),
    .D1(_10631_),
    .Y(_10646_));
 sky130_fd_sc_hd__a22o_1 _20856_ (.A1(_10631_),
    .A2(_10633_),
    .B1(_10639_),
    .B2(_10643_),
    .X(_10647_));
 sky130_fd_sc_hd__o22ai_4 _20857_ (.A1(_12670_),
    .A2(net327),
    .B1(_10634_),
    .B2(_10644_),
    .Y(_10648_));
 sky130_fd_sc_hd__o211ai_2 _20858_ (.A1(_12670_),
    .A2(net327),
    .B1(_10646_),
    .C1(_10647_),
    .Y(_10649_));
 sky130_fd_sc_hd__o22ai_4 _20859_ (.A1(net311),
    .A2(_10626_),
    .B1(_10645_),
    .B2(_10648_),
    .Y(_10650_));
 sky130_fd_sc_hd__inv_2 _20860_ (.A(_10650_),
    .Y(_10652_));
 sky130_fd_sc_hd__and3_1 _20861_ (.A(_00022_),
    .B(_00044_),
    .C(_10650_),
    .X(_10653_));
 sky130_fd_sc_hd__a211o_2 _20862_ (.A1(_10628_),
    .A2(_10649_),
    .B1(_00011_),
    .C1(net323),
    .X(_10654_));
 sky130_fd_sc_hd__a311oi_4 _20863_ (.A1(_10647_),
    .A2(net311),
    .A3(_10646_),
    .B1(net232),
    .C1(_10627_),
    .Y(_10655_));
 sky130_fd_sc_hd__o221ai_4 _20864_ (.A1(net311),
    .A2(_10626_),
    .B1(_10645_),
    .B2(_10648_),
    .C1(net234),
    .Y(_10656_));
 sky130_fd_sc_hd__a2bb2oi_1 _20865_ (.A1_N(_06622_),
    .A2_N(_06624_),
    .B1(_10628_),
    .B2(_10649_),
    .Y(_10657_));
 sky130_fd_sc_hd__o21ai_4 _20866_ (.A1(_06622_),
    .A2(_06624_),
    .B1(_10650_),
    .Y(_10658_));
 sky130_fd_sc_hd__a21oi_1 _20867_ (.A1(_09758_),
    .A2(_10192_),
    .B1(_10194_),
    .Y(_10659_));
 sky130_fd_sc_hd__a31o_1 _20868_ (.A1(_09761_),
    .A2(_10191_),
    .A3(_10195_),
    .B1(_10196_),
    .X(_10660_));
 sky130_fd_sc_hd__a21oi_1 _20869_ (.A1(_10193_),
    .A2(_10195_),
    .B1(_10196_),
    .Y(_10661_));
 sky130_fd_sc_hd__a21oi_2 _20870_ (.A1(_10656_),
    .A2(_10658_),
    .B1(_10660_),
    .Y(_10663_));
 sky130_fd_sc_hd__o21bai_4 _20871_ (.A1(_10655_),
    .A2(_10657_),
    .B1_N(_10660_),
    .Y(_10664_));
 sky130_fd_sc_hd__o2bb2ai_1 _20872_ (.A1_N(net232),
    .A2_N(_10650_),
    .B1(_10659_),
    .B2(_10196_),
    .Y(_10665_));
 sky130_fd_sc_hd__nand3_4 _20873_ (.A(_10656_),
    .B(_10658_),
    .C(_10660_),
    .Y(_10666_));
 sky130_fd_sc_hd__o22ai_4 _20874_ (.A1(_00011_),
    .A2(net323),
    .B1(_10655_),
    .B2(_10665_),
    .Y(_10667_));
 sky130_fd_sc_hd__nand3_2 _20875_ (.A(_10664_),
    .B(_10666_),
    .C(net307),
    .Y(_10668_));
 sky130_fd_sc_hd__o22ai_4 _20876_ (.A1(net308),
    .A2(_10652_),
    .B1(_10663_),
    .B2(_10667_),
    .Y(_10669_));
 sky130_fd_sc_hd__o221a_1 _20877_ (.A1(net262),
    .A2(_09775_),
    .B1(net254),
    .B2(_10206_),
    .C1(_10213_),
    .X(_10670_));
 sky130_fd_sc_hd__a31oi_4 _20878_ (.A1(_09778_),
    .A2(_10207_),
    .A3(_10213_),
    .B1(_10208_),
    .Y(_10671_));
 sky130_fd_sc_hd__a31oi_2 _20879_ (.A1(_10664_),
    .A2(_10666_),
    .A3(net307),
    .B1(net251),
    .Y(_10672_));
 sky130_fd_sc_hd__a311oi_4 _20880_ (.A1(_10664_),
    .A2(_10666_),
    .A3(net308),
    .B1(net251),
    .C1(_10653_),
    .Y(_10674_));
 sky130_fd_sc_hd__o221ai_4 _20881_ (.A1(net308),
    .A2(_10652_),
    .B1(_10663_),
    .B2(_10667_),
    .C1(_06314_),
    .Y(_10675_));
 sky130_fd_sc_hd__a2bb2oi_4 _20882_ (.A1_N(_06305_),
    .A2_N(_06307_),
    .B1(_10654_),
    .B2(_10668_),
    .Y(_10676_));
 sky130_fd_sc_hd__o21ai_1 _20883_ (.A1(_06305_),
    .A2(_06307_),
    .B1(_10669_),
    .Y(_10677_));
 sky130_fd_sc_hd__a21oi_1 _20884_ (.A1(_10654_),
    .A2(_10672_),
    .B1(_10676_),
    .Y(_10678_));
 sky130_fd_sc_hd__o211ai_1 _20885_ (.A1(_10208_),
    .A2(_10670_),
    .B1(_10675_),
    .C1(_10677_),
    .Y(_10679_));
 sky130_fd_sc_hd__o21ai_1 _20886_ (.A1(_10674_),
    .A2(_10676_),
    .B1(_10671_),
    .Y(_10680_));
 sky130_fd_sc_hd__nand3_2 _20887_ (.A(_10679_),
    .B(_10680_),
    .C(net279),
    .Y(_10681_));
 sky130_fd_sc_hd__a21oi_2 _20888_ (.A1(_10654_),
    .A2(_10668_),
    .B1(net279),
    .Y(_10682_));
 sky130_fd_sc_hd__a211o_1 _20889_ (.A1(_10654_),
    .A2(_10668_),
    .B1(_01940_),
    .C1(_01951_),
    .X(_10683_));
 sky130_fd_sc_hd__nand3_2 _20890_ (.A(_10677_),
    .B(_10671_),
    .C(_10675_),
    .Y(_10685_));
 sky130_fd_sc_hd__o22ai_4 _20891_ (.A1(_10208_),
    .A2(_10670_),
    .B1(_10674_),
    .B2(_10676_),
    .Y(_10686_));
 sky130_fd_sc_hd__o211ai_4 _20892_ (.A1(_01940_),
    .A2(_01951_),
    .B1(_10685_),
    .C1(_10686_),
    .Y(_10687_));
 sky130_fd_sc_hd__a31o_2 _20893_ (.A1(_10685_),
    .A2(_10686_),
    .A3(net279),
    .B1(_10682_),
    .X(_10688_));
 sky130_fd_sc_hd__a31oi_4 _20894_ (.A1(_10685_),
    .A2(_10686_),
    .A3(net279),
    .B1(_10682_),
    .Y(_10689_));
 sky130_fd_sc_hd__a2bb2oi_1 _20895_ (.A1_N(_06009_),
    .A2_N(_06010_),
    .B1(_10683_),
    .B2(_10687_),
    .Y(_10690_));
 sky130_fd_sc_hd__o211ai_4 _20896_ (.A1(_10669_),
    .A2(net279),
    .B1(net253),
    .C1(_10681_),
    .Y(_10691_));
 sky130_fd_sc_hd__o211a_1 _20897_ (.A1(net286),
    .A2(_06012_),
    .B1(_10683_),
    .C1(_10687_),
    .X(_10692_));
 sky130_fd_sc_hd__o211ai_4 _20898_ (.A1(net286),
    .A2(_06012_),
    .B1(_10683_),
    .C1(_10687_),
    .Y(_10693_));
 sky130_fd_sc_hd__nand2_1 _20899_ (.A(_10691_),
    .B(_10693_),
    .Y(_10694_));
 sky130_fd_sc_hd__a22o_1 _20900_ (.A1(net261),
    .A2(_10217_),
    .B1(_10224_),
    .B2(_10226_),
    .X(_10696_));
 sky130_fd_sc_hd__a31oi_4 _20901_ (.A1(_10220_),
    .A2(_10224_),
    .A3(_10226_),
    .B1(_10218_),
    .Y(_10697_));
 sky130_fd_sc_hd__a22oi_4 _20902_ (.A1(_10691_),
    .A2(_10693_),
    .B1(_10696_),
    .B2(_10220_),
    .Y(_10698_));
 sky130_fd_sc_hd__nand4_2 _20903_ (.A(_10219_),
    .B(_10228_),
    .C(_10691_),
    .D(_10693_),
    .Y(_10699_));
 sky130_fd_sc_hd__o2bb2ai_1 _20904_ (.A1_N(_10219_),
    .A2_N(_10228_),
    .B1(_10690_),
    .B2(_10692_),
    .Y(_10700_));
 sky130_fd_sc_hd__o211ai_4 _20905_ (.A1(net302),
    .A2(_04019_),
    .B1(_10699_),
    .C1(_10700_),
    .Y(_10701_));
 sky130_fd_sc_hd__o211a_1 _20906_ (.A1(_10669_),
    .A2(net279),
    .B1(_04040_),
    .C1(_10681_),
    .X(_10702_));
 sky130_fd_sc_hd__o22ai_4 _20907_ (.A1(_04008_),
    .A2(_04019_),
    .B1(_10697_),
    .B2(_10694_),
    .Y(_10703_));
 sky130_fd_sc_hd__a2bb2o_2 _20908_ (.A1_N(_10703_),
    .A2_N(_10698_),
    .B1(_10688_),
    .B2(_04040_),
    .X(_10704_));
 sky130_fd_sc_hd__o22a_4 _20909_ (.A1(net276),
    .A2(_10689_),
    .B1(_10698_),
    .B2(_10703_),
    .X(_10705_));
 sky130_fd_sc_hd__nand4_2 _20910_ (.A(_08950_),
    .B(_08953_),
    .C(_09361_),
    .D(_09362_),
    .Y(_10707_));
 sky130_fd_sc_hd__a211oi_4 _20911_ (.A1(_09800_),
    .A2(_09821_),
    .B1(_10707_),
    .C1(_09824_),
    .Y(_10708_));
 sky130_fd_sc_hd__nand2_1 _20912_ (.A(_10240_),
    .B(_10708_),
    .Y(_10709_));
 sky130_fd_sc_hd__o211ai_4 _20913_ (.A1(_10244_),
    .A2(_10239_),
    .B1(_10242_),
    .C1(_10709_),
    .Y(_10710_));
 sky130_fd_sc_hd__o211ai_4 _20914_ (.A1(net267),
    .A2(_10235_),
    .B1(_10708_),
    .C1(_08956_),
    .Y(_10711_));
 sky130_fd_sc_hd__nand4_4 _20915_ (.A(_10708_),
    .B(_10242_),
    .C(_10240_),
    .D(_08956_),
    .Y(_10712_));
 sky130_fd_sc_hd__o21ai_4 _20916_ (.A1(_10239_),
    .A2(_10711_),
    .B1(_10710_),
    .Y(_10713_));
 sky130_fd_sc_hd__o211a_1 _20917_ (.A1(net276),
    .A2(_10688_),
    .B1(_10701_),
    .C1(net261),
    .X(_10714_));
 sky130_fd_sc_hd__o211ai_4 _20918_ (.A1(net276),
    .A2(_10688_),
    .B1(_10701_),
    .C1(net261),
    .Y(_10715_));
 sky130_fd_sc_hd__o22ai_2 _20919_ (.A1(_05765_),
    .A2(net289),
    .B1(_10698_),
    .B2(_10703_),
    .Y(_10716_));
 sky130_fd_sc_hd__o221a_1 _20920_ (.A1(net276),
    .A2(_10689_),
    .B1(_10698_),
    .B2(_10703_),
    .C1(net262),
    .X(_10718_));
 sky130_fd_sc_hd__o221ai_4 _20921_ (.A1(net276),
    .A2(_10689_),
    .B1(_10698_),
    .B2(_10703_),
    .C1(net262),
    .Y(_10719_));
 sky130_fd_sc_hd__o21a_1 _20922_ (.A1(_10702_),
    .A2(_10716_),
    .B1(_10715_),
    .X(_10720_));
 sky130_fd_sc_hd__o21ai_1 _20923_ (.A1(_10702_),
    .A2(_10716_),
    .B1(_10715_),
    .Y(_10721_));
 sky130_fd_sc_hd__a21oi_2 _20924_ (.A1(_10710_),
    .A2(_10712_),
    .B1(_10721_),
    .Y(_10722_));
 sky130_fd_sc_hd__o22ai_2 _20925_ (.A1(net297),
    .A2(_05232_),
    .B1(_10720_),
    .B2(_10713_),
    .Y(_10723_));
 sky130_fd_sc_hd__o2bb2ai_1 _20926_ (.A1_N(_10710_),
    .A2_N(_10712_),
    .B1(_10714_),
    .B2(_10718_),
    .Y(_10724_));
 sky130_fd_sc_hd__nand4_1 _20927_ (.A(_10710_),
    .B(_10712_),
    .C(_10715_),
    .D(_10719_),
    .Y(_10725_));
 sky130_fd_sc_hd__o221a_1 _20928_ (.A1(_05228_),
    .A2(_05230_),
    .B1(_10688_),
    .B2(net276),
    .C1(_10701_),
    .X(_10726_));
 sky130_fd_sc_hd__nand3_2 _20929_ (.A(_10724_),
    .B(_10725_),
    .C(net273),
    .Y(_10727_));
 sky130_fd_sc_hd__a31o_2 _20930_ (.A1(_10724_),
    .A2(_10725_),
    .A3(net273),
    .B1(_10726_),
    .X(_10729_));
 sky130_fd_sc_hd__inv_2 _20931_ (.A(_10729_),
    .Y(_10730_));
 sky130_fd_sc_hd__o221a_2 _20932_ (.A1(net273),
    .A2(_10704_),
    .B1(_10722_),
    .B2(_10723_),
    .C1(_05486_),
    .X(_10731_));
 sky130_fd_sc_hd__o21ai_2 _20933_ (.A1(_05478_),
    .A2(_05479_),
    .B1(_10729_),
    .Y(_10732_));
 sky130_fd_sc_hd__o311a_1 _20934_ (.A1(net297),
    .A2(_05232_),
    .A3(_10705_),
    .B1(net267),
    .C1(_10727_),
    .X(_10733_));
 sky130_fd_sc_hd__o211ai_4 _20935_ (.A1(net273),
    .A2(_10705_),
    .B1(net267),
    .C1(_10727_),
    .Y(_10734_));
 sky130_fd_sc_hd__o221ai_4 _20936_ (.A1(net273),
    .A2(_10704_),
    .B1(_10722_),
    .B2(_10723_),
    .C1(net291),
    .Y(_10735_));
 sky130_fd_sc_hd__a21oi_1 _20937_ (.A1(net294),
    .A2(_10252_),
    .B1(_10257_),
    .Y(_10736_));
 sky130_fd_sc_hd__o21ai_1 _20938_ (.A1(_09835_),
    .A2(_10255_),
    .B1(_10259_),
    .Y(_10737_));
 sky130_fd_sc_hd__a21o_1 _20939_ (.A1(_10259_),
    .A2(_10257_),
    .B1(_10260_),
    .X(_10738_));
 sky130_fd_sc_hd__a21oi_1 _20940_ (.A1(_10259_),
    .A2(_10257_),
    .B1(_10260_),
    .Y(_10740_));
 sky130_fd_sc_hd__o2bb2ai_2 _20941_ (.A1_N(_10734_),
    .A2_N(_10735_),
    .B1(_10736_),
    .B2(_10258_),
    .Y(_10741_));
 sky130_fd_sc_hd__a22oi_2 _20942_ (.A1(_10261_),
    .A2(_10737_),
    .B1(_10729_),
    .B2(net292),
    .Y(_10742_));
 sky130_fd_sc_hd__nand3_2 _20943_ (.A(_10738_),
    .B(_10735_),
    .C(_10734_),
    .Y(_10743_));
 sky130_fd_sc_hd__nand3_2 _20944_ (.A(_10741_),
    .B(_10743_),
    .C(net246),
    .Y(_10744_));
 sky130_fd_sc_hd__a31o_1 _20945_ (.A1(_10741_),
    .A2(_10743_),
    .A3(net246),
    .B1(_10731_),
    .X(_10745_));
 sky130_fd_sc_hd__o22a_1 _20946_ (.A1(_09852_),
    .A2(_10275_),
    .B1(net299),
    .B2(_10270_),
    .X(_10746_));
 sky130_fd_sc_hd__nand2_1 _20947_ (.A(_10274_),
    .B(_10276_),
    .Y(_10747_));
 sky130_fd_sc_hd__o21ai_2 _20948_ (.A1(net299),
    .A2(_10270_),
    .B1(_10747_),
    .Y(_10748_));
 sky130_fd_sc_hd__a311oi_4 _20949_ (.A1(_10741_),
    .A2(_10743_),
    .A3(net246),
    .B1(_10731_),
    .C1(net294),
    .Y(_10749_));
 sky130_fd_sc_hd__a311o_1 _20950_ (.A1(_10741_),
    .A2(_10743_),
    .A3(net246),
    .B1(_10731_),
    .C1(net294),
    .X(_10751_));
 sky130_fd_sc_hd__a2bb2oi_2 _20951_ (.A1_N(net318),
    .A2_N(_05244_),
    .B1(_10732_),
    .B2(_10744_),
    .Y(_10752_));
 sky130_fd_sc_hd__a22o_1 _20952_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_10732_),
    .B2(_10744_),
    .X(_10753_));
 sky130_fd_sc_hd__o211ai_1 _20953_ (.A1(_10273_),
    .A2(_10746_),
    .B1(_10751_),
    .C1(_10753_),
    .Y(_10754_));
 sky130_fd_sc_hd__o2bb2ai_1 _20954_ (.A1_N(_10272_),
    .A2_N(_10747_),
    .B1(_10749_),
    .B2(_10752_),
    .Y(_10755_));
 sky130_fd_sc_hd__nand3_1 _20955_ (.A(_10754_),
    .B(_10755_),
    .C(net242),
    .Y(_10756_));
 sky130_fd_sc_hd__a21oi_2 _20956_ (.A1(_10732_),
    .A2(_10744_),
    .B1(net242),
    .Y(_10757_));
 sky130_fd_sc_hd__a211o_1 _20957_ (.A1(_10732_),
    .A2(_10744_),
    .B1(net266),
    .C1(_05751_),
    .X(_10758_));
 sky130_fd_sc_hd__nand3_2 _20958_ (.A(_10753_),
    .B(_10748_),
    .C(_10751_),
    .Y(_10759_));
 sky130_fd_sc_hd__o22ai_4 _20959_ (.A1(_10273_),
    .A2(_10746_),
    .B1(_10749_),
    .B2(_10752_),
    .Y(_10760_));
 sky130_fd_sc_hd__nand3_1 _20960_ (.A(_10759_),
    .B(_10760_),
    .C(net242),
    .Y(_10762_));
 sky130_fd_sc_hd__a31oi_4 _20961_ (.A1(_10759_),
    .A2(_10760_),
    .A3(net242),
    .B1(_10757_),
    .Y(_10763_));
 sky130_fd_sc_hd__o211a_1 _20962_ (.A1(_10745_),
    .A2(net242),
    .B1(net298),
    .C1(_10756_),
    .X(_10764_));
 sky130_fd_sc_hd__o211ai_4 _20963_ (.A1(_10745_),
    .A2(net242),
    .B1(net298),
    .C1(_10756_),
    .Y(_10765_));
 sky130_fd_sc_hd__a311oi_4 _20964_ (.A1(_10759_),
    .A2(_10760_),
    .A3(net242),
    .B1(_10757_),
    .C1(net298),
    .Y(_10766_));
 sky130_fd_sc_hd__o211ai_2 _20965_ (.A1(_04206_),
    .A2(_04216_),
    .B1(_10758_),
    .C1(_10762_),
    .Y(_10767_));
 sky130_fd_sc_hd__a21oi_1 _20966_ (.A1(_10302_),
    .A2(_10305_),
    .B1(_10290_),
    .Y(_10768_));
 sky130_fd_sc_hd__a31o_1 _20967_ (.A1(_10294_),
    .A2(_10302_),
    .A3(_10305_),
    .B1(_10290_),
    .X(_10769_));
 sky130_fd_sc_hd__o2bb2ai_2 _20968_ (.A1_N(_10765_),
    .A2_N(_10767_),
    .B1(_10768_),
    .B2(_10293_),
    .Y(_10770_));
 sky130_fd_sc_hd__o2bb2ai_1 _20969_ (.A1_N(_10291_),
    .A2_N(_10315_),
    .B1(net299),
    .B2(_10763_),
    .Y(_10771_));
 sky130_fd_sc_hd__a31oi_1 _20970_ (.A1(_10769_),
    .A2(_10767_),
    .A3(_10765_),
    .B1(_05995_),
    .Y(_10773_));
 sky130_fd_sc_hd__o221ai_4 _20971_ (.A1(net259),
    .A2(net257),
    .B1(_10766_),
    .B2(_10771_),
    .C1(_10770_),
    .Y(_10774_));
 sky130_fd_sc_hd__or3_4 _20972_ (.A(net259),
    .B(net257),
    .C(_10763_),
    .X(_10775_));
 sky130_fd_sc_hd__a2bb2o_1 _20973_ (.A1_N(net240),
    .A2_N(_10763_),
    .B1(_10770_),
    .B2(_10773_),
    .X(_10776_));
 sky130_fd_sc_hd__a21oi_4 _20974_ (.A1(_10774_),
    .A2(_10775_),
    .B1(_02137_),
    .Y(_10777_));
 sky130_fd_sc_hd__a22o_1 _20975_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_10774_),
    .B2(_10775_),
    .X(_10778_));
 sky130_fd_sc_hd__a21oi_1 _20976_ (.A1(_10773_),
    .A2(_10770_),
    .B1(_02148_),
    .Y(_10779_));
 sky130_fd_sc_hd__o311a_1 _20977_ (.A1(net259),
    .A2(net257),
    .A3(_10763_),
    .B1(_02137_),
    .C1(_10774_),
    .X(_10780_));
 sky130_fd_sc_hd__o211ai_4 _20978_ (.A1(net240),
    .A2(_10763_),
    .B1(_02137_),
    .C1(_10774_),
    .Y(_10781_));
 sky130_fd_sc_hd__nand4_1 _20979_ (.A(_09016_),
    .B(_09019_),
    .C(_09431_),
    .D(_09433_),
    .Y(_10782_));
 sky130_fd_sc_hd__nor3_1 _20980_ (.A(_10782_),
    .B(_09891_),
    .C(_09889_),
    .Y(_10784_));
 sky130_fd_sc_hd__nand3b_1 _20981_ (.A_N(_10782_),
    .B(_09892_),
    .C(_09890_),
    .Y(_10785_));
 sky130_fd_sc_hd__a31oi_1 _20982_ (.A1(_10317_),
    .A2(_00240_),
    .A3(_10313_),
    .B1(_10785_),
    .Y(_10786_));
 sky130_fd_sc_hd__a31o_1 _20983_ (.A1(_10317_),
    .A2(_00240_),
    .A3(_10313_),
    .B1(_10785_),
    .X(_10787_));
 sky130_fd_sc_hd__a32oi_1 _20984_ (.A1(_00251_),
    .A2(_10288_),
    .A3(_10310_),
    .B1(_10324_),
    .B2(_10784_),
    .Y(_10788_));
 sky130_fd_sc_hd__a211oi_2 _20985_ (.A1(_10328_),
    .A2(_10324_),
    .B1(_10325_),
    .C1(_10786_),
    .Y(_10789_));
 sky130_fd_sc_hd__o211ai_4 _20986_ (.A1(_10329_),
    .A2(_10323_),
    .B1(_10326_),
    .C1(_10787_),
    .Y(_10790_));
 sky130_fd_sc_hd__nand3_2 _20987_ (.A(_10324_),
    .B(_10784_),
    .C(_09022_),
    .Y(_10791_));
 sky130_fd_sc_hd__and3_1 _20988_ (.A(_09022_),
    .B(_10786_),
    .C(_10326_),
    .X(_10792_));
 sky130_fd_sc_hd__nand4_1 _20989_ (.A(_10324_),
    .B(_10326_),
    .C(_10784_),
    .D(_09022_),
    .Y(_10793_));
 sky130_fd_sc_hd__a2bb2oi_2 _20990_ (.A1_N(_10325_),
    .A2_N(_10791_),
    .B1(_10332_),
    .B2(_10788_),
    .Y(_10795_));
 sky130_fd_sc_hd__o21ai_1 _20991_ (.A1(_10325_),
    .A2(_10791_),
    .B1(_10781_),
    .Y(_10796_));
 sky130_fd_sc_hd__o2111ai_4 _20992_ (.A1(_10791_),
    .A2(_10325_),
    .B1(_10781_),
    .C1(_10790_),
    .D1(_10778_),
    .Y(_10797_));
 sky130_fd_sc_hd__a21oi_2 _20993_ (.A1(_10775_),
    .A2(_10779_),
    .B1(_10777_),
    .Y(_10798_));
 sky130_fd_sc_hd__o22ai_4 _20994_ (.A1(_10777_),
    .A2(_10780_),
    .B1(_10789_),
    .B2(_10792_),
    .Y(_10799_));
 sky130_fd_sc_hd__o211ai_4 _20995_ (.A1(_10795_),
    .A2(_10798_),
    .B1(_10797_),
    .C1(net212),
    .Y(_10800_));
 sky130_fd_sc_hd__a21oi_4 _20996_ (.A1(_10774_),
    .A2(_10775_),
    .B1(net213),
    .Y(_10801_));
 sky130_fd_sc_hd__a22o_2 _20997_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_10774_),
    .B2(_10775_),
    .X(_10802_));
 sky130_fd_sc_hd__a31oi_4 _20998_ (.A1(_10799_),
    .A2(net213),
    .A3(_10797_),
    .B1(_10801_),
    .Y(_10803_));
 sky130_fd_sc_hd__a21oi_4 _20999_ (.A1(_10800_),
    .A2(_10802_),
    .B1(net211),
    .Y(_10804_));
 sky130_fd_sc_hd__or3_1 _21000_ (.A(_06608_),
    .B(net237),
    .C(_10803_),
    .X(_10806_));
 sky130_fd_sc_hd__a31o_1 _21001_ (.A1(_10799_),
    .A2(net213),
    .A3(_10797_),
    .B1(_00251_),
    .X(_10807_));
 sky130_fd_sc_hd__a311oi_4 _21002_ (.A1(_10799_),
    .A2(net213),
    .A3(_10797_),
    .B1(_10801_),
    .C1(_00251_),
    .Y(_10808_));
 sky130_fd_sc_hd__nand3_2 _21003_ (.A(_10800_),
    .B(_10802_),
    .C(_00240_),
    .Y(_10809_));
 sky130_fd_sc_hd__a21oi_1 _21004_ (.A1(_10800_),
    .A2(_10802_),
    .B1(_00240_),
    .Y(_10810_));
 sky130_fd_sc_hd__a21o_2 _21005_ (.A1(_10800_),
    .A2(_10802_),
    .B1(_00240_),
    .X(_10811_));
 sky130_fd_sc_hd__o32a_1 _21006_ (.A1(net361),
    .A2(net345),
    .A3(_10336_),
    .B1(_10339_),
    .B2(_10342_),
    .X(_10812_));
 sky130_fd_sc_hd__a21oi_2 _21007_ (.A1(_10341_),
    .A2(_10339_),
    .B1(_10342_),
    .Y(_10813_));
 sky130_fd_sc_hd__o21ai_4 _21008_ (.A1(_10808_),
    .A2(_10810_),
    .B1(_10813_),
    .Y(_10814_));
 sky130_fd_sc_hd__o211ai_4 _21009_ (.A1(_10801_),
    .A2(_10807_),
    .B1(_10812_),
    .C1(_10811_),
    .Y(_10815_));
 sky130_fd_sc_hd__nand3_1 _21010_ (.A(_10814_),
    .B(_10815_),
    .C(net211),
    .Y(_10817_));
 sky130_fd_sc_hd__a31oi_4 _21011_ (.A1(_10814_),
    .A2(_10815_),
    .A3(net211),
    .B1(_10804_),
    .Y(_10818_));
 sky130_fd_sc_hd__a31o_1 _21012_ (.A1(_10814_),
    .A2(_10815_),
    .A3(net211),
    .B1(_10804_),
    .X(_10819_));
 sky130_fd_sc_hd__o311a_1 _21013_ (.A1(net365),
    .A2(net364),
    .A3(_09917_),
    .B1(_09925_),
    .C1(_10353_),
    .X(_10820_));
 sky130_fd_sc_hd__a21bo_1 _21014_ (.A1(_10354_),
    .A2(_10358_),
    .B1_N(_10353_),
    .X(_10821_));
 sky130_fd_sc_hd__a311oi_4 _21015_ (.A1(_10814_),
    .A2(_10815_),
    .A3(net211),
    .B1(_10804_),
    .C1(net326),
    .Y(_10822_));
 sky130_fd_sc_hd__o221ai_2 _21016_ (.A1(_12867_),
    .A2(_12877_),
    .B1(net211),
    .B2(_10803_),
    .C1(_10817_),
    .Y(_10823_));
 sky130_fd_sc_hd__a2bb2oi_1 _21017_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_10806_),
    .B2(_10817_),
    .Y(_10824_));
 sky130_fd_sc_hd__a2bb2o_1 _21018_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_10806_),
    .B2(_10817_),
    .X(_10825_));
 sky130_fd_sc_hd__o211ai_1 _21019_ (.A1(_10356_),
    .A2(_10820_),
    .B1(_10823_),
    .C1(_10825_),
    .Y(_10826_));
 sky130_fd_sc_hd__o21ai_1 _21020_ (.A1(_10822_),
    .A2(_10824_),
    .B1(_10821_),
    .Y(_10828_));
 sky130_fd_sc_hd__nand3_1 _21021_ (.A(_10826_),
    .B(_10828_),
    .C(net208),
    .Y(_10829_));
 sky130_fd_sc_hd__and3_1 _21022_ (.A(_06900_),
    .B(_06902_),
    .C(_10819_),
    .X(_10830_));
 sky130_fd_sc_hd__or3_1 _21023_ (.A(net230),
    .B(_06901_),
    .C(_10818_),
    .X(_10831_));
 sky130_fd_sc_hd__o21ai_2 _21024_ (.A1(_12888_),
    .A2(_10818_),
    .B1(_10821_),
    .Y(_10832_));
 sky130_fd_sc_hd__o22ai_2 _21025_ (.A1(_10356_),
    .A2(_10820_),
    .B1(_10822_),
    .B2(_10824_),
    .Y(_10833_));
 sky130_fd_sc_hd__o221a_1 _21026_ (.A1(net230),
    .A2(_06901_),
    .B1(_10822_),
    .B2(_10832_),
    .C1(_10833_),
    .X(_10834_));
 sky130_fd_sc_hd__o221ai_4 _21027_ (.A1(net230),
    .A2(_06901_),
    .B1(_10822_),
    .B2(_10832_),
    .C1(_10833_),
    .Y(_10835_));
 sky130_fd_sc_hd__a31o_1 _21028_ (.A1(_06900_),
    .A2(_06902_),
    .A3(_10819_),
    .B1(_10834_),
    .X(_10836_));
 sky130_fd_sc_hd__o31a_2 _21029_ (.A1(net230),
    .A2(_06901_),
    .A3(_10818_),
    .B1(_10835_),
    .X(_10837_));
 sky130_fd_sc_hd__a2bb2oi_2 _21030_ (.A1_N(_11210_),
    .A2_N(_11232_),
    .B1(_10831_),
    .B2(_10835_),
    .Y(_10839_));
 sky130_fd_sc_hd__o211ai_4 _21031_ (.A1(_10819_),
    .A2(net208),
    .B1(_11309_),
    .C1(_10829_),
    .Y(_10840_));
 sky130_fd_sc_hd__o211a_1 _21032_ (.A1(net208),
    .A2(_10818_),
    .B1(_11298_),
    .C1(_10835_),
    .X(_10841_));
 sky130_fd_sc_hd__o211ai_4 _21033_ (.A1(net208),
    .A2(_10818_),
    .B1(_11298_),
    .C1(_10835_),
    .Y(_10842_));
 sky130_fd_sc_hd__a21o_1 _21034_ (.A1(_10370_),
    .A2(_10371_),
    .B1(_10367_),
    .X(_10843_));
 sky130_fd_sc_hd__o2111ai_1 _21035_ (.A1(_10015_),
    .A2(_10365_),
    .B1(_10374_),
    .C1(_10840_),
    .D1(_10842_),
    .Y(_10844_));
 sky130_fd_sc_hd__o22ai_1 _21036_ (.A1(_10367_),
    .A2(_10373_),
    .B1(_10839_),
    .B2(_10841_),
    .Y(_10845_));
 sky130_fd_sc_hd__o211ai_2 _21037_ (.A1(_07227_),
    .A2(net203),
    .B1(_10844_),
    .C1(_10845_),
    .Y(_10846_));
 sky130_fd_sc_hd__a21oi_2 _21038_ (.A1(_10840_),
    .A2(_10842_),
    .B1(_10843_),
    .Y(_10847_));
 sky130_fd_sc_hd__a31o_1 _21039_ (.A1(_10840_),
    .A2(_10842_),
    .A3(_10843_),
    .B1(_07232_),
    .X(_10848_));
 sky130_fd_sc_hd__o22ai_4 _21040_ (.A1(net185),
    .A2(_10837_),
    .B1(_10847_),
    .B2(_10848_),
    .Y(_10850_));
 sky130_fd_sc_hd__o211ai_4 _21041_ (.A1(_10836_),
    .A2(net185),
    .B1(_10025_),
    .C1(_10846_),
    .Y(_10851_));
 sky130_fd_sc_hd__o221ai_4 _21042_ (.A1(net185),
    .A2(_10837_),
    .B1(_10847_),
    .B2(_10848_),
    .C1(_10015_),
    .Y(_10852_));
 sky130_fd_sc_hd__inv_2 _21043_ (.A(_10852_),
    .Y(_10853_));
 sky130_fd_sc_hd__o22a_2 _21044_ (.A1(_09953_),
    .A2(_09955_),
    .B1(_08918_),
    .B2(_10381_),
    .X(_10854_));
 sky130_fd_sc_hd__o21ai_1 _21045_ (.A1(_10383_),
    .A2(_10384_),
    .B1(_10387_),
    .Y(_10855_));
 sky130_fd_sc_hd__o2bb2ai_1 _21046_ (.A1_N(_10851_),
    .A2_N(_10852_),
    .B1(_10854_),
    .B2(_10386_),
    .Y(_10856_));
 sky130_fd_sc_hd__o2111ai_4 _21047_ (.A1(_10383_),
    .A2(_10384_),
    .B1(_10387_),
    .C1(_10851_),
    .D1(_10852_),
    .Y(_10857_));
 sky130_fd_sc_hd__a21o_1 _21048_ (.A1(_10851_),
    .A2(_10852_),
    .B1(_10855_),
    .X(_10858_));
 sky130_fd_sc_hd__o21ai_2 _21049_ (.A1(_10386_),
    .A2(_10854_),
    .B1(_10852_),
    .Y(_10859_));
 sky130_fd_sc_hd__o221ai_4 _21050_ (.A1(_10386_),
    .A2(_10854_),
    .B1(_10025_),
    .B2(_10850_),
    .C1(_10851_),
    .Y(_10861_));
 sky130_fd_sc_hd__a22oi_4 _21051_ (.A1(_07545_),
    .A2(_07547_),
    .B1(_10856_),
    .B2(_10857_),
    .Y(_10862_));
 sky130_fd_sc_hd__nand3_2 _21052_ (.A(_10858_),
    .B(_10861_),
    .C(net163),
    .Y(_10863_));
 sky130_fd_sc_hd__o311a_1 _21053_ (.A1(net185),
    .A2(_10830_),
    .A3(_10834_),
    .B1(_10846_),
    .C1(_07550_),
    .X(_10864_));
 sky130_fd_sc_hd__nand2_1 _21054_ (.A(_10850_),
    .B(_07550_),
    .Y(_10865_));
 sky130_fd_sc_hd__a21oi_4 _21055_ (.A1(_07550_),
    .A2(_10850_),
    .B1(_10862_),
    .Y(_10866_));
 sky130_fd_sc_hd__or3_2 _21056_ (.A(_07912_),
    .B(_07914_),
    .C(_10866_),
    .X(_10867_));
 sky130_fd_sc_hd__o21ai_1 _21057_ (.A1(_10405_),
    .A2(_10401_),
    .B1(_10400_),
    .Y(_10868_));
 sky130_fd_sc_hd__a311oi_1 _21058_ (.A1(_10858_),
    .A2(_10861_),
    .A3(net163),
    .B1(_10864_),
    .C1(_08918_),
    .Y(_10869_));
 sky130_fd_sc_hd__o211ai_2 _21059_ (.A1(_08863_),
    .A2(_08885_),
    .B1(_10863_),
    .C1(_10865_),
    .Y(_10870_));
 sky130_fd_sc_hd__a21oi_4 _21060_ (.A1(_10863_),
    .A2(_10865_),
    .B1(_08907_),
    .Y(_10872_));
 sky130_fd_sc_hd__o22ai_1 _21061_ (.A1(_08819_),
    .A2(_08841_),
    .B1(_10862_),
    .B2(_10864_),
    .Y(_10873_));
 sky130_fd_sc_hd__o211ai_2 _21062_ (.A1(_10398_),
    .A2(_10409_),
    .B1(_10870_),
    .C1(_10873_),
    .Y(_10874_));
 sky130_fd_sc_hd__o21bai_1 _21063_ (.A1(_10869_),
    .A2(_10872_),
    .B1_N(_10868_),
    .Y(_10875_));
 sky130_fd_sc_hd__nand3_4 _21064_ (.A(_10875_),
    .B(net160),
    .C(_10874_),
    .Y(_10876_));
 sky130_fd_sc_hd__o21ai_4 _21065_ (.A1(net160),
    .A2(_10866_),
    .B1(_10876_),
    .Y(_10877_));
 sky130_fd_sc_hd__o221a_1 _21066_ (.A1(_09977_),
    .A2(_09978_),
    .B1(_10415_),
    .B2(_07033_),
    .C1(_09975_),
    .X(_10878_));
 sky130_fd_sc_hd__o32a_1 _21067_ (.A1(_06945_),
    .A2(_06967_),
    .A3(_10416_),
    .B1(_09981_),
    .B2(_09974_),
    .X(_10879_));
 sky130_fd_sc_hd__o32a_1 _21068_ (.A1(_06945_),
    .A2(_06967_),
    .A3(_10416_),
    .B1(_10019_),
    .B2(_10419_),
    .X(_10880_));
 sky130_fd_sc_hd__o221a_2 _21069_ (.A1(net368),
    .A2(_07866_),
    .B1(net160),
    .B2(_10866_),
    .C1(_10876_),
    .X(_10881_));
 sky130_fd_sc_hd__o221ai_4 _21070_ (.A1(net368),
    .A2(_07866_),
    .B1(net160),
    .B2(_10866_),
    .C1(_10876_),
    .Y(_10883_));
 sky130_fd_sc_hd__a21oi_4 _21071_ (.A1(_10867_),
    .A2(_10876_),
    .B1(_07888_),
    .Y(_10884_));
 sky130_fd_sc_hd__a22o_1 _21072_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_10867_),
    .B2(_10876_),
    .X(_10885_));
 sky130_fd_sc_hd__o211ai_1 _21073_ (.A1(_10417_),
    .A2(_10878_),
    .B1(_10883_),
    .C1(_10885_),
    .Y(_10886_));
 sky130_fd_sc_hd__o22ai_1 _21074_ (.A1(_10419_),
    .A2(_10879_),
    .B1(_10881_),
    .B2(_10884_),
    .Y(_10887_));
 sky130_fd_sc_hd__nand3_1 _21075_ (.A(_10886_),
    .B(_10887_),
    .C(_08300_),
    .Y(_10888_));
 sky130_fd_sc_hd__a211o_1 _21076_ (.A1(_10867_),
    .A2(_10876_),
    .B1(net180),
    .C1(_08298_),
    .X(_10889_));
 sky130_fd_sc_hd__o22a_1 _21077_ (.A1(_10419_),
    .A2(_10879_),
    .B1(_10877_),
    .B2(_07899_),
    .X(_10890_));
 sky130_fd_sc_hd__o21ai_2 _21078_ (.A1(_10419_),
    .A2(_10879_),
    .B1(_10883_),
    .Y(_10891_));
 sky130_fd_sc_hd__o22ai_1 _21079_ (.A1(_10417_),
    .A2(_10878_),
    .B1(_10881_),
    .B2(_10884_),
    .Y(_10892_));
 sky130_fd_sc_hd__o211ai_2 _21080_ (.A1(_10884_),
    .A2(_10891_),
    .B1(_08300_),
    .C1(_10892_),
    .Y(_10894_));
 sky130_fd_sc_hd__o21ai_2 _21081_ (.A1(_08300_),
    .A2(_10877_),
    .B1(_10888_),
    .Y(_10895_));
 sky130_fd_sc_hd__o211ai_4 _21082_ (.A1(_06989_),
    .A2(net375),
    .B1(_10889_),
    .C1(_10894_),
    .Y(_10896_));
 sky130_fd_sc_hd__inv_2 _21083_ (.A(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__a2bb2oi_1 _21084_ (.A1_N(_06945_),
    .A2_N(_06967_),
    .B1(_10889_),
    .B2(_10894_),
    .Y(_10898_));
 sky130_fd_sc_hd__o211ai_2 _21085_ (.A1(_10877_),
    .A2(_08300_),
    .B1(_07044_),
    .C1(_10888_),
    .Y(_10899_));
 sky130_fd_sc_hd__nand3_1 _21086_ (.A(_10484_),
    .B(_10896_),
    .C(_10899_),
    .Y(_10900_));
 sky130_fd_sc_hd__a21o_1 _21087_ (.A1(_10896_),
    .A2(_10899_),
    .B1(_10484_),
    .X(_10901_));
 sky130_fd_sc_hd__o211ai_4 _21088_ (.A1(net158),
    .A2(_08712_),
    .B1(_10900_),
    .C1(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__or3_2 _21089_ (.A(net158),
    .B(_08712_),
    .C(_10895_),
    .X(_10903_));
 sky130_fd_sc_hd__o21ai_1 _21090_ (.A1(_08714_),
    .A2(_10895_),
    .B1(_10902_),
    .Y(_10905_));
 sky130_fd_sc_hd__a21oi_4 _21091_ (.A1(_10902_),
    .A2(_10903_),
    .B1(_06332_),
    .Y(_10906_));
 sky130_fd_sc_hd__o221a_1 _21092_ (.A1(net381),
    .A2(_06310_),
    .B1(_08714_),
    .B2(_10895_),
    .C1(_10902_),
    .X(_10907_));
 sky130_fd_sc_hd__o221ai_2 _21093_ (.A1(net381),
    .A2(_06310_),
    .B1(_08714_),
    .B2(_10895_),
    .C1(_10902_),
    .Y(_10908_));
 sky130_fd_sc_hd__a31o_1 _21094_ (.A1(_10429_),
    .A2(_10439_),
    .A3(_10446_),
    .B1(_10445_),
    .X(_10909_));
 sky130_fd_sc_hd__a31oi_4 _21095_ (.A1(_10429_),
    .A2(_10439_),
    .A3(_10446_),
    .B1(_10445_),
    .Y(_10910_));
 sky130_fd_sc_hd__o21ai_1 _21096_ (.A1(_10906_),
    .A2(_10907_),
    .B1(_10910_),
    .Y(_10911_));
 sky130_fd_sc_hd__o21ai_1 _21097_ (.A1(_10906_),
    .A2(_10907_),
    .B1(_10909_),
    .Y(_10912_));
 sky130_fd_sc_hd__o21a_1 _21098_ (.A1(_06343_),
    .A2(_10905_),
    .B1(_10910_),
    .X(_10913_));
 sky130_fd_sc_hd__a31o_1 _21099_ (.A1(_10902_),
    .A2(_10903_),
    .A3(_06332_),
    .B1(_10909_),
    .X(_10914_));
 sky130_fd_sc_hd__o311ai_2 _21100_ (.A1(_10906_),
    .A2(_10910_),
    .A3(_10907_),
    .B1(_09125_),
    .C1(_10911_),
    .Y(_10916_));
 sky130_fd_sc_hd__o221ai_4 _21101_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_10906_),
    .B2(_10914_),
    .C1(_10912_),
    .Y(_10917_));
 sky130_fd_sc_hd__a211o_1 _21102_ (.A1(_10902_),
    .A2(_10903_),
    .B1(_09120_),
    .C1(_09121_),
    .X(_10918_));
 sky130_fd_sc_hd__o311ai_2 _21103_ (.A1(_10448_),
    .A2(_10441_),
    .A3(_10440_),
    .B1(_10455_),
    .C1(_10450_),
    .Y(_10919_));
 sky130_fd_sc_hd__nand2_1 _21104_ (.A(_10456_),
    .B(_10919_),
    .Y(_10920_));
 sky130_fd_sc_hd__a22o_1 _21105_ (.A1(net395),
    .A2(_05796_),
    .B1(_10456_),
    .B2(_10919_),
    .X(_10921_));
 sky130_fd_sc_hd__and3_1 _21106_ (.A(_10919_),
    .B(_05851_),
    .C(_10456_),
    .X(_10922_));
 sky130_fd_sc_hd__o221a_1 _21107_ (.A1(_09553_),
    .A2(net155),
    .B1(_10920_),
    .B2(_05862_),
    .C1(_10921_),
    .X(_10923_));
 sky130_fd_sc_hd__o221ai_2 _21108_ (.A1(_05862_),
    .A2(_10920_),
    .B1(net155),
    .B2(_09553_),
    .C1(_10921_),
    .Y(_10924_));
 sky130_fd_sc_hd__o211ai_2 _21109_ (.A1(_09125_),
    .A2(_10905_),
    .B1(_10923_),
    .C1(_10916_),
    .Y(_10925_));
 sky130_fd_sc_hd__nand3_2 _21110_ (.A(_10917_),
    .B(_10918_),
    .C(_10924_),
    .Y(_10927_));
 sky130_fd_sc_hd__nand2_1 _21111_ (.A(_10925_),
    .B(_10927_),
    .Y(_10928_));
 sky130_fd_sc_hd__o21ai_1 _21112_ (.A1(_10013_),
    .A2(_10462_),
    .B1(_10463_),
    .Y(_10929_));
 sky130_fd_sc_hd__o221ai_4 _21113_ (.A1(_05501_),
    .A2(_05523_),
    .B1(_10013_),
    .B2(_10462_),
    .C1(_10463_),
    .Y(_10930_));
 sky130_fd_sc_hd__o21ai_2 _21114_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_10929_),
    .Y(_10931_));
 sky130_fd_sc_hd__o211ai_2 _21115_ (.A1(_09571_),
    .A2(_09573_),
    .B1(_10930_),
    .C1(_10931_),
    .Y(_10932_));
 sky130_fd_sc_hd__a21o_1 _21116_ (.A1(_10925_),
    .A2(_10927_),
    .B1(_10932_),
    .X(_10933_));
 sky130_fd_sc_hd__a31o_1 _21117_ (.A1(_09579_),
    .A2(_10930_),
    .A3(_10931_),
    .B1(_10928_),
    .X(_10934_));
 sky130_fd_sc_hd__nand3b_1 _21118_ (.A_N(_10932_),
    .B(_10927_),
    .C(_10925_),
    .Y(_10935_));
 sky130_fd_sc_hd__nand2_1 _21119_ (.A(_10928_),
    .B(_10932_),
    .Y(_10936_));
 sky130_fd_sc_hd__nand2_1 _21120_ (.A(_10933_),
    .B(_10934_),
    .Y(_10938_));
 sky130_fd_sc_hd__a21o_1 _21121_ (.A1(_10933_),
    .A2(_10934_),
    .B1(_05250_),
    .X(_10939_));
 sky130_fd_sc_hd__a21oi_1 _21122_ (.A1(_10935_),
    .A2(_10936_),
    .B1(_05239_),
    .Y(_10940_));
 sky130_fd_sc_hd__a21o_1 _21123_ (.A1(_10935_),
    .A2(_10936_),
    .B1(_05239_),
    .X(_10941_));
 sky130_fd_sc_hd__a21oi_1 _21124_ (.A1(_10939_),
    .A2(_10941_),
    .B1(_10470_),
    .Y(_10942_));
 sky130_fd_sc_hd__a31o_1 _21125_ (.A1(_10939_),
    .A2(_10941_),
    .A3(_10470_),
    .B1(_10479_),
    .X(_10943_));
 sky130_fd_sc_hd__a2bb2o_1 _21126_ (.A1_N(_10942_),
    .A2_N(_10943_),
    .B1(_10479_),
    .B2(_10938_),
    .X(_10944_));
 sky130_fd_sc_hd__nand2_1 _21127_ (.A(_10944_),
    .B(net1),
    .Y(_10945_));
 sky130_fd_sc_hd__xor2_1 _21128_ (.A(net1),
    .B(_10944_),
    .X(_10946_));
 sky130_fd_sc_hd__or4_4 _21129_ (.A(net51),
    .B(net52),
    .C(net53),
    .D(_09552_),
    .X(_10947_));
 sky130_fd_sc_hd__and3b_4 _21130_ (.A_N(net54),
    .B(_10947_),
    .C(net57),
    .X(_10949_));
 sky130_fd_sc_hd__inv_6 _21131_ (.A(net137),
    .Y(_10950_));
 sky130_fd_sc_hd__a21boi_4 _21132_ (.A1(_10947_),
    .A2(net57),
    .B1_N(net54),
    .Y(_10951_));
 sky130_fd_sc_hd__a21bo_4 _21133_ (.A1(_10947_),
    .A2(net57),
    .B1_N(net54),
    .X(_10952_));
 sky130_fd_sc_hd__nor2_8 _21134_ (.A(_10949_),
    .B(net136),
    .Y(_10953_));
 sky130_fd_sc_hd__nand2_8 _21135_ (.A(_10950_),
    .B(_10952_),
    .Y(_10954_));
 sky130_fd_sc_hd__or3_1 _21136_ (.A(_10949_),
    .B(net136),
    .C(_10944_),
    .X(_10955_));
 sky130_fd_sc_hd__o21ai_2 _21137_ (.A1(_10946_),
    .A2(_10953_),
    .B1(_10955_),
    .Y(_10956_));
 sky130_fd_sc_hd__o21ai_1 _21138_ (.A1(_05051_),
    .A2(_10483_),
    .B1(_10956_),
    .Y(_10957_));
 sky130_fd_sc_hd__or3_1 _21139_ (.A(_05051_),
    .B(_10483_),
    .C(_10956_),
    .X(_10958_));
 sky130_fd_sc_hd__and2_1 _21140_ (.A(_10957_),
    .B(_10958_),
    .X(net86));
 sky130_fd_sc_hd__o2bb2a_1 _21141_ (.A1_N(_10483_),
    .A2_N(_10956_),
    .B1(_04832_),
    .B2(_04942_),
    .X(_10960_));
 sky130_fd_sc_hd__a21oi_2 _21142_ (.A1(_10908_),
    .A2(_10910_),
    .B1(_10906_),
    .Y(_10961_));
 sky130_fd_sc_hd__or4_4 _21143_ (.A(net20),
    .B(net21),
    .C(net22),
    .D(_09586_),
    .X(_10962_));
 sky130_fd_sc_hd__or3b_4 _21144_ (.A(_03399_),
    .B(net24),
    .C_N(_10962_),
    .X(_10963_));
 sky130_fd_sc_hd__a21bo_4 _21145_ (.A1(_10962_),
    .A2(net410),
    .B1_N(net24),
    .X(_10964_));
 sky130_fd_sc_hd__o311a_4 _21146_ (.A1(net21),
    .A2(net22),
    .A3(_10020_),
    .B1(net24),
    .C1(net410),
    .X(_10965_));
 sky130_fd_sc_hd__o211ai_4 _21147_ (.A1(net22),
    .A2(_10485_),
    .B1(net24),
    .C1(net410),
    .Y(_10966_));
 sky130_fd_sc_hd__a21oi_4 _21148_ (.A1(_10962_),
    .A2(net410),
    .B1(net24),
    .Y(_10967_));
 sky130_fd_sc_hd__a21o_4 _21149_ (.A1(_10962_),
    .A2(net410),
    .B1(net24),
    .X(_10968_));
 sky130_fd_sc_hd__nand2_8 _21150_ (.A(_10966_),
    .B(_10968_),
    .Y(_10970_));
 sky130_fd_sc_hd__nor2_8 _21151_ (.A(_10965_),
    .B(_10967_),
    .Y(_10971_));
 sky130_fd_sc_hd__a31o_1 _21152_ (.A1(_10968_),
    .A2(net33),
    .A3(_10966_),
    .B1(net405),
    .X(_10972_));
 sky130_fd_sc_hd__o32a_1 _21153_ (.A1(_03178_),
    .A2(_10965_),
    .A3(_10967_),
    .B1(_10489_),
    .B2(_10490_),
    .X(_10973_));
 sky130_fd_sc_hd__and3_1 _21154_ (.A(_10971_),
    .B(net33),
    .C(_10492_),
    .X(_10974_));
 sky130_fd_sc_hd__or4_1 _21155_ (.A(_03178_),
    .B(_10489_),
    .C(_10490_),
    .D(_10970_),
    .X(_10975_));
 sky130_fd_sc_hd__or2_1 _21156_ (.A(_10973_),
    .B(_10974_),
    .X(_10976_));
 sky130_fd_sc_hd__o221a_1 _21157_ (.A1(_10029_),
    .A2(net150),
    .B1(_10973_),
    .B2(_10974_),
    .C1(_10505_),
    .X(_10977_));
 sky130_fd_sc_hd__o221ai_2 _21158_ (.A1(_10029_),
    .A2(net150),
    .B1(_10973_),
    .B2(_10974_),
    .C1(_10505_),
    .Y(_10978_));
 sky130_fd_sc_hd__a21oi_2 _21159_ (.A1(_10501_),
    .A2(_10505_),
    .B1(_10976_),
    .Y(_10979_));
 sky130_fd_sc_hd__a21o_1 _21160_ (.A1(_10501_),
    .A2(_10505_),
    .B1(_10976_),
    .X(_10981_));
 sky130_fd_sc_hd__o21ai_1 _21161_ (.A1(_10977_),
    .A2(_10979_),
    .B1(net405),
    .Y(_10982_));
 sky130_fd_sc_hd__and3_1 _21162_ (.A(_10971_),
    .B(net33),
    .C(_05185_),
    .X(_10983_));
 sky130_fd_sc_hd__or4_1 _21163_ (.A(_03178_),
    .B(net405),
    .C(_10965_),
    .D(_10967_),
    .X(_10984_));
 sky130_fd_sc_hd__o31a_1 _21164_ (.A1(_05185_),
    .A2(_10977_),
    .A3(_10979_),
    .B1(_10984_),
    .X(_10985_));
 sky130_fd_sc_hd__or3_2 _21165_ (.A(_05348_),
    .B(net401),
    .C(_10985_),
    .X(_10986_));
 sky130_fd_sc_hd__and3_1 _21166_ (.A(net151),
    .B(_10972_),
    .C(_10982_),
    .X(_10987_));
 sky130_fd_sc_hd__o211ai_1 _21167_ (.A1(_10021_),
    .A2(_10022_),
    .B1(_10972_),
    .C1(_10982_),
    .Y(_10988_));
 sky130_fd_sc_hd__o311a_1 _21168_ (.A1(_05185_),
    .A2(_10977_),
    .A3(_10979_),
    .B1(_10984_),
    .C1(net153),
    .X(_10989_));
 sky130_fd_sc_hd__a311o_1 _21169_ (.A1(_10981_),
    .A2(net405),
    .A3(_10978_),
    .B1(_10983_),
    .C1(net151),
    .X(_10990_));
 sky130_fd_sc_hd__o211ai_1 _21170_ (.A1(_10023_),
    .A2(_10024_),
    .B1(_10972_),
    .C1(_10982_),
    .Y(_10992_));
 sky130_fd_sc_hd__a311o_1 _21171_ (.A1(_10981_),
    .A2(net405),
    .A3(_10978_),
    .B1(_10983_),
    .C1(net153),
    .X(_10993_));
 sky130_fd_sc_hd__nand2_1 _21172_ (.A(_10992_),
    .B(_10993_),
    .Y(_10994_));
 sky130_fd_sc_hd__nand2_1 _21173_ (.A(_10988_),
    .B(_10990_),
    .Y(_10995_));
 sky130_fd_sc_hd__nand4_2 _21174_ (.A(_10044_),
    .B(_09160_),
    .C(_10043_),
    .D(_09611_),
    .Y(_10996_));
 sky130_fd_sc_hd__a21oi_1 _21175_ (.A1(_09163_),
    .A2(_09166_),
    .B1(_10996_),
    .Y(_10997_));
 sky130_fd_sc_hd__nor4_2 _21176_ (.A(_09167_),
    .B(_10512_),
    .C(_10996_),
    .D(_10515_),
    .Y(_10998_));
 sky130_fd_sc_hd__nand2_1 _21177_ (.A(_10517_),
    .B(_10997_),
    .Y(_10999_));
 sky130_fd_sc_hd__o2bb2a_1 _21178_ (.A1_N(_10507_),
    .A2_N(_10514_),
    .B1(_10512_),
    .B2(_10996_),
    .X(_11000_));
 sky130_fd_sc_hd__o21ai_1 _21179_ (.A1(_10512_),
    .A2(_10996_),
    .B1(_10516_),
    .Y(_11001_));
 sky130_fd_sc_hd__a31oi_2 _21180_ (.A1(_10517_),
    .A2(_10518_),
    .A3(_10043_),
    .B1(_11001_),
    .Y(_11003_));
 sky130_fd_sc_hd__a31o_1 _21181_ (.A1(_10517_),
    .A2(_10518_),
    .A3(_10043_),
    .B1(_11001_),
    .X(_11004_));
 sky130_fd_sc_hd__o22ai_2 _21182_ (.A1(_10987_),
    .A2(_10989_),
    .B1(_10998_),
    .B2(_11003_),
    .Y(_11005_));
 sky130_fd_sc_hd__a211oi_2 _21183_ (.A1(_10520_),
    .A2(_11000_),
    .B1(_10998_),
    .C1(_10995_),
    .Y(_11006_));
 sky130_fd_sc_hd__nand3_4 _21184_ (.A(_11004_),
    .B(_10994_),
    .C(_10999_),
    .Y(_11007_));
 sky130_fd_sc_hd__nand3_2 _21185_ (.A(_05403_),
    .B(_11005_),
    .C(_11007_),
    .Y(_11008_));
 sky130_fd_sc_hd__o311a_1 _21186_ (.A1(_05185_),
    .A2(_10977_),
    .A3(_10979_),
    .B1(_10984_),
    .C1(_05392_),
    .X(_11009_));
 sky130_fd_sc_hd__a21oi_2 _21187_ (.A1(_11005_),
    .A2(_11007_),
    .B1(_05392_),
    .Y(_11010_));
 sky130_fd_sc_hd__o31a_1 _21188_ (.A1(_05348_),
    .A2(net401),
    .A3(_10985_),
    .B1(_11008_),
    .X(_11011_));
 sky130_fd_sc_hd__o21ai_1 _21189_ (.A1(_05403_),
    .A2(_10985_),
    .B1(_11008_),
    .Y(_11012_));
 sky130_fd_sc_hd__or4_2 _21190_ (.A(_05676_),
    .B(_05698_),
    .C(_11009_),
    .D(_11010_),
    .X(_11014_));
 sky130_fd_sc_hd__o221ai_4 _21191_ (.A1(net177),
    .A2(_10054_),
    .B1(_10523_),
    .B2(net174),
    .C1(_10067_),
    .Y(_11015_));
 sky130_fd_sc_hd__a31oi_1 _21192_ (.A1(_05403_),
    .A2(_11005_),
    .A3(_11007_),
    .B1(_09595_),
    .Y(_11016_));
 sky130_fd_sc_hd__o211a_1 _21193_ (.A1(_05403_),
    .A2(_10985_),
    .B1(net172),
    .C1(_11008_),
    .X(_11017_));
 sky130_fd_sc_hd__nand3_1 _21194_ (.A(_11008_),
    .B(net172),
    .C(_10986_),
    .Y(_11018_));
 sky130_fd_sc_hd__a2bb2oi_2 _21195_ (.A1_N(_09588_),
    .A2_N(net187),
    .B1(_10986_),
    .B2(_11008_),
    .Y(_11019_));
 sky130_fd_sc_hd__a21oi_2 _21196_ (.A1(_10986_),
    .A2(_11016_),
    .B1(_11019_),
    .Y(_11020_));
 sky130_fd_sc_hd__o211ai_2 _21197_ (.A1(net173),
    .A2(_10524_),
    .B1(_11015_),
    .C1(_11020_),
    .Y(_11021_));
 sky130_fd_sc_hd__o22ai_2 _21198_ (.A1(net174),
    .A2(_10523_),
    .B1(_11017_),
    .B2(_11019_),
    .Y(_11022_));
 sky130_fd_sc_hd__o211ai_4 _21199_ (.A1(_10531_),
    .A2(_11022_),
    .B1(_11021_),
    .C1(net358),
    .Y(_11023_));
 sky130_fd_sc_hd__o21ai_1 _21200_ (.A1(net358),
    .A2(_11011_),
    .B1(_11023_),
    .Y(_11025_));
 sky130_fd_sc_hd__o311a_2 _21201_ (.A1(net358),
    .A2(_11009_),
    .A3(_11010_),
    .B1(_11023_),
    .C1(_06848_),
    .X(_11026_));
 sky130_fd_sc_hd__o32ai_1 _21202_ (.A1(net177),
    .A2(_10525_),
    .A3(_10535_),
    .B1(_10547_),
    .B2(_10548_),
    .Y(_11027_));
 sky130_fd_sc_hd__a2bb2oi_2 _21203_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_11014_),
    .B2(_11023_),
    .Y(_11028_));
 sky130_fd_sc_hd__a2bb2o_2 _21204_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_11014_),
    .B2(_11023_),
    .X(_11029_));
 sky130_fd_sc_hd__o211a_1 _21205_ (.A1(net358),
    .A2(_11011_),
    .B1(net174),
    .C1(_11023_),
    .X(_11030_));
 sky130_fd_sc_hd__o211ai_2 _21206_ (.A1(net358),
    .A2(_11011_),
    .B1(net174),
    .C1(_11023_),
    .Y(_11031_));
 sky130_fd_sc_hd__nor2_1 _21207_ (.A(_11028_),
    .B(_11030_),
    .Y(_11032_));
 sky130_fd_sc_hd__nand2_2 _21208_ (.A(_11027_),
    .B(_11032_),
    .Y(_11033_));
 sky130_fd_sc_hd__o221ai_4 _21209_ (.A1(_11028_),
    .A2(_11030_),
    .B1(_10547_),
    .B2(_10548_),
    .C1(_10543_),
    .Y(_11034_));
 sky130_fd_sc_hd__a22oi_4 _21210_ (.A1(_06804_),
    .A2(_06826_),
    .B1(_11033_),
    .B2(_11034_),
    .Y(_11036_));
 sky130_fd_sc_hd__a211o_2 _21211_ (.A1(_11014_),
    .A2(_11023_),
    .B1(_06793_),
    .C1(_06815_),
    .X(_11037_));
 sky130_fd_sc_hd__nand3_4 _21212_ (.A(_11033_),
    .B(_11034_),
    .C(net357),
    .Y(_11038_));
 sky130_fd_sc_hd__a31o_2 _21213_ (.A1(_06848_),
    .A2(_11014_),
    .A3(_11023_),
    .B1(_11036_),
    .X(_11039_));
 sky130_fd_sc_hd__a21oi_2 _21214_ (.A1(_11037_),
    .A2(_11038_),
    .B1(net355),
    .Y(_11040_));
 sky130_fd_sc_hd__or4_1 _21215_ (.A(net374),
    .B(_07702_),
    .C(_11026_),
    .D(_11036_),
    .X(_11041_));
 sky130_fd_sc_hd__a2bb2oi_1 _21216_ (.A1_N(_08724_),
    .A2_N(_08726_),
    .B1(_11037_),
    .B2(_11038_),
    .Y(_11042_));
 sky130_fd_sc_hd__a22o_2 _21217_ (.A1(_08725_),
    .A2(_08727_),
    .B1(_11037_),
    .B2(_11038_),
    .X(_11043_));
 sky130_fd_sc_hd__and3_1 _21218_ (.A(_11038_),
    .B(net177),
    .C(_11037_),
    .X(_11044_));
 sky130_fd_sc_hd__o211ai_4 _21219_ (.A1(_08728_),
    .A2(net195),
    .B1(_11037_),
    .C1(_11038_),
    .Y(_11045_));
 sky130_fd_sc_hd__o41ai_4 _21220_ (.A1(_08728_),
    .A2(net195),
    .A3(_11026_),
    .A4(_11036_),
    .B1(_11045_),
    .Y(_11047_));
 sky130_fd_sc_hd__a22oi_4 _21221_ (.A1(net198),
    .A2(_10557_),
    .B1(_10575_),
    .B2(_10566_),
    .Y(_11048_));
 sky130_fd_sc_hd__o221ai_4 _21222_ (.A1(net199),
    .A2(_10556_),
    .B1(_11042_),
    .B2(_11044_),
    .C1(_10578_),
    .Y(_11049_));
 sky130_fd_sc_hd__o221a_1 _21223_ (.A1(net374),
    .A2(_07702_),
    .B1(_11047_),
    .B2(_11048_),
    .C1(_11049_),
    .X(_11050_));
 sky130_fd_sc_hd__o221ai_4 _21224_ (.A1(net374),
    .A2(_07702_),
    .B1(_11047_),
    .B2(_11048_),
    .C1(_11049_),
    .Y(_11051_));
 sky130_fd_sc_hd__o31a_4 _21225_ (.A1(net354),
    .A2(_11026_),
    .A3(_11036_),
    .B1(_11051_),
    .X(_11052_));
 sky130_fd_sc_hd__inv_2 _21226_ (.A(_11052_),
    .Y(_11053_));
 sky130_fd_sc_hd__a2bb2oi_1 _21227_ (.A1_N(_08307_),
    .A2_N(_08309_),
    .B1(_11041_),
    .B2(_11051_),
    .Y(_11054_));
 sky130_fd_sc_hd__o22ai_4 _21228_ (.A1(_08307_),
    .A2(_08309_),
    .B1(_11040_),
    .B2(_11050_),
    .Y(_11055_));
 sky130_fd_sc_hd__o221a_1 _21229_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_11039_),
    .B2(net354),
    .C1(_11051_),
    .X(_11056_));
 sky130_fd_sc_hd__o221ai_4 _21230_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_11039_),
    .B2(net354),
    .C1(_11051_),
    .Y(_11058_));
 sky130_fd_sc_hd__nor2_1 _21231_ (.A(_11054_),
    .B(_11056_),
    .Y(_11059_));
 sky130_fd_sc_hd__nand2_1 _21232_ (.A(_11055_),
    .B(_11058_),
    .Y(_11060_));
 sky130_fd_sc_hd__nor3b_2 _21233_ (.A(_09689_),
    .B(_09691_),
    .C_N(_09232_),
    .Y(_11061_));
 sky130_fd_sc_hd__and3_1 _21234_ (.A(_11061_),
    .B(_10125_),
    .C(_10121_),
    .X(_11062_));
 sky130_fd_sc_hd__and4_1 _21235_ (.A(_11061_),
    .B(_10125_),
    .C(_10121_),
    .D(_09241_),
    .X(_11063_));
 sky130_fd_sc_hd__nand4_1 _21236_ (.A(_11061_),
    .B(_10125_),
    .C(_10121_),
    .D(_09241_),
    .Y(_11064_));
 sky130_fd_sc_hd__nand3_1 _21237_ (.A(_10590_),
    .B(_11061_),
    .C(_10126_),
    .Y(_11065_));
 sky130_fd_sc_hd__nand4_4 _21238_ (.A(_11062_),
    .B(_10592_),
    .C(_10590_),
    .D(_09241_),
    .Y(_11066_));
 sky130_fd_sc_hd__a31oi_1 _21239_ (.A1(_10126_),
    .A2(_10590_),
    .A3(_11061_),
    .B1(_10591_),
    .Y(_11067_));
 sky130_fd_sc_hd__o211a_1 _21240_ (.A1(_10589_),
    .A2(_10588_),
    .B1(_11065_),
    .C1(_10592_),
    .X(_11069_));
 sky130_fd_sc_hd__o211ai_4 _21241_ (.A1(_10589_),
    .A2(_10588_),
    .B1(_11065_),
    .C1(_10592_),
    .Y(_11070_));
 sky130_fd_sc_hd__a22oi_2 _21242_ (.A1(_10593_),
    .A2(_11063_),
    .B1(_11067_),
    .B2(_10594_),
    .Y(_11071_));
 sky130_fd_sc_hd__a31o_1 _21243_ (.A1(_09241_),
    .A2(_10593_),
    .A3(_11062_),
    .B1(_11069_),
    .X(_11072_));
 sky130_fd_sc_hd__a21oi_1 _21244_ (.A1(_11066_),
    .A2(_11070_),
    .B1(_11060_),
    .Y(_11073_));
 sky130_fd_sc_hd__o211ai_1 _21245_ (.A1(_11054_),
    .A2(_11056_),
    .B1(_11066_),
    .C1(_11070_),
    .Y(_11074_));
 sky130_fd_sc_hd__o21ai_1 _21246_ (.A1(_08678_),
    .A2(_08700_),
    .B1(_11074_),
    .Y(_11075_));
 sky130_fd_sc_hd__nand4_4 _21247_ (.A(_11055_),
    .B(_11058_),
    .C(_11066_),
    .D(_11070_),
    .Y(_11076_));
 sky130_fd_sc_hd__a22o_1 _21248_ (.A1(_11055_),
    .A2(_11058_),
    .B1(_11066_),
    .B2(_11070_),
    .X(_11077_));
 sky130_fd_sc_hd__o221ai_4 _21249_ (.A1(_08678_),
    .A2(_08700_),
    .B1(_11059_),
    .B2(_11071_),
    .C1(_11076_),
    .Y(_11078_));
 sky130_fd_sc_hd__o211a_1 _21250_ (.A1(_11040_),
    .A2(_11050_),
    .B1(_08689_),
    .C1(_08711_),
    .X(_11080_));
 sky130_fd_sc_hd__or3_1 _21251_ (.A(_08678_),
    .B(_08700_),
    .C(_11052_),
    .X(_11081_));
 sky130_fd_sc_hd__a31o_1 _21252_ (.A1(_11077_),
    .A2(net338),
    .A3(_11076_),
    .B1(_11080_),
    .X(_11082_));
 sky130_fd_sc_hd__a211o_2 _21253_ (.A1(_11078_),
    .A2(_11081_),
    .B1(net351),
    .C1(_09807_),
    .X(_11083_));
 sky130_fd_sc_hd__o211a_1 _21254_ (.A1(net224),
    .A2(_10136_),
    .B1(_10144_),
    .C1(_10600_),
    .X(_11084_));
 sky130_fd_sc_hd__a22o_1 _21255_ (.A1(net202),
    .A2(_10598_),
    .B1(_10604_),
    .B2(_10140_),
    .X(_11085_));
 sky130_fd_sc_hd__o211a_1 _21256_ (.A1(net222),
    .A2(_10134_),
    .B1(_10602_),
    .C1(_10604_),
    .X(_11086_));
 sky130_fd_sc_hd__a22oi_2 _21257_ (.A1(_07929_),
    .A2(_07932_),
    .B1(_11078_),
    .B2(_11081_),
    .Y(_11087_));
 sky130_fd_sc_hd__o221ai_4 _21258_ (.A1(net338),
    .A2(_11053_),
    .B1(_11073_),
    .B2(_11075_),
    .C1(_07936_),
    .Y(_11088_));
 sky130_fd_sc_hd__a311oi_4 _21259_ (.A1(_11077_),
    .A2(net338),
    .A3(_11076_),
    .B1(_11080_),
    .C1(_07936_),
    .Y(_11089_));
 sky130_fd_sc_hd__o211ai_4 _21260_ (.A1(net338),
    .A2(_11052_),
    .B1(_07935_),
    .C1(_11078_),
    .Y(_11091_));
 sky130_fd_sc_hd__o21ai_1 _21261_ (.A1(_10599_),
    .A2(_11086_),
    .B1(_11091_),
    .Y(_11092_));
 sky130_fd_sc_hd__o211a_1 _21262_ (.A1(_10599_),
    .A2(_11086_),
    .B1(_11088_),
    .C1(_11091_),
    .X(_11093_));
 sky130_fd_sc_hd__o2111ai_4 _21263_ (.A1(net202),
    .A2(_10598_),
    .B1(_11085_),
    .C1(_11088_),
    .D1(_11091_),
    .Y(_11094_));
 sky130_fd_sc_hd__a22oi_2 _21264_ (.A1(_10602_),
    .A2(_11085_),
    .B1(_11088_),
    .B2(_11091_),
    .Y(_11095_));
 sky130_fd_sc_hd__o22ai_2 _21265_ (.A1(_10601_),
    .A2(_11084_),
    .B1(_11087_),
    .B2(_11089_),
    .Y(_11096_));
 sky130_fd_sc_hd__nand3_2 _21266_ (.A(_11096_),
    .B(net335),
    .C(_11094_),
    .Y(_11097_));
 sky130_fd_sc_hd__o21ai_1 _21267_ (.A1(_11093_),
    .A2(_11095_),
    .B1(net335),
    .Y(_11098_));
 sky130_fd_sc_hd__o31a_2 _21268_ (.A1(_09840_),
    .A2(_11093_),
    .A3(_11095_),
    .B1(_11083_),
    .X(_11099_));
 sky130_fd_sc_hd__inv_2 _21269_ (.A(_11099_),
    .Y(_11100_));
 sky130_fd_sc_hd__a2bb2oi_4 _21270_ (.A1_N(_07555_),
    .A2_N(net218),
    .B1(_11083_),
    .B2(_11097_),
    .Y(_11102_));
 sky130_fd_sc_hd__o221ai_4 _21271_ (.A1(_07555_),
    .A2(net218),
    .B1(_11082_),
    .B2(net335),
    .C1(_11098_),
    .Y(_11103_));
 sky130_fd_sc_hd__a31oi_1 _21272_ (.A1(_11096_),
    .A2(net335),
    .A3(_11094_),
    .B1(net202),
    .Y(_11104_));
 sky130_fd_sc_hd__o311a_1 _21273_ (.A1(_09840_),
    .A2(_11093_),
    .A3(_11095_),
    .B1(_07564_),
    .C1(_11083_),
    .X(_11105_));
 sky130_fd_sc_hd__nand3_4 _21274_ (.A(_11097_),
    .B(_07564_),
    .C(_11083_),
    .Y(_11106_));
 sky130_fd_sc_hd__a21oi_2 _21275_ (.A1(_11083_),
    .A2(_11104_),
    .B1(_11102_),
    .Y(_11107_));
 sky130_fd_sc_hd__o211ai_4 _21276_ (.A1(net227),
    .A2(_10149_),
    .B1(_10615_),
    .C1(_10620_),
    .Y(_11108_));
 sky130_fd_sc_hd__o2bb2ai_2 _21277_ (.A1_N(_10152_),
    .A2_N(_10620_),
    .B1(_10613_),
    .B2(net222),
    .Y(_11109_));
 sky130_fd_sc_hd__o21ai_2 _21278_ (.A1(net222),
    .A2(_10613_),
    .B1(_11108_),
    .Y(_11110_));
 sky130_fd_sc_hd__o2111ai_4 _21279_ (.A1(_10614_),
    .A2(net224),
    .B1(_11106_),
    .C1(_11103_),
    .D1(_11109_),
    .Y(_11111_));
 sky130_fd_sc_hd__o221ai_4 _21280_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_11110_),
    .B2(_11107_),
    .C1(_11111_),
    .Y(_11113_));
 sky130_fd_sc_hd__or3_1 _21281_ (.A(_11046_),
    .B(_11057_),
    .C(_11099_),
    .X(_11114_));
 sky130_fd_sc_hd__o21ai_1 _21282_ (.A1(_11102_),
    .A2(_11105_),
    .B1(_11110_),
    .Y(_11115_));
 sky130_fd_sc_hd__o2111ai_4 _21283_ (.A1(_10613_),
    .A2(net222),
    .B1(_11106_),
    .C1(_11103_),
    .D1(_11108_),
    .Y(_11116_));
 sky130_fd_sc_hd__nand3_4 _21284_ (.A(_11115_),
    .B(_11116_),
    .C(net332),
    .Y(_11117_));
 sky130_fd_sc_hd__o21ai_4 _21285_ (.A1(net332),
    .A2(_11099_),
    .B1(_11117_),
    .Y(_11118_));
 sky130_fd_sc_hd__inv_2 _21286_ (.A(_11118_),
    .Y(_11119_));
 sky130_fd_sc_hd__o211ai_4 _21287_ (.A1(_11100_),
    .A2(net332),
    .B1(net222),
    .C1(_11113_),
    .Y(_11120_));
 sky130_fd_sc_hd__and3_1 _21288_ (.A(_11117_),
    .B(net224),
    .C(_11114_),
    .X(_11121_));
 sky130_fd_sc_hd__o211ai_4 _21289_ (.A1(net332),
    .A2(_11099_),
    .B1(net224),
    .C1(_11117_),
    .Y(_11122_));
 sky130_fd_sc_hd__nand2_1 _21290_ (.A(_11120_),
    .B(_11122_),
    .Y(_11124_));
 sky130_fd_sc_hd__o211ai_2 _21291_ (.A1(_10641_),
    .A2(_08886_),
    .B1(_10633_),
    .C1(_10639_),
    .Y(_11125_));
 sky130_fd_sc_hd__a31oi_2 _21292_ (.A1(_10633_),
    .A2(_10639_),
    .A3(_10643_),
    .B1(_10630_),
    .Y(_11126_));
 sky130_fd_sc_hd__o311a_2 _21293_ (.A1(_06918_),
    .A2(_06920_),
    .A3(_10626_),
    .B1(_10646_),
    .C1(_11124_),
    .X(_11127_));
 sky130_fd_sc_hd__o211ai_2 _21294_ (.A1(net227),
    .A2(_10626_),
    .B1(_10646_),
    .C1(_11124_),
    .Y(_11128_));
 sky130_fd_sc_hd__o2111ai_4 _21295_ (.A1(_10630_),
    .A2(_10644_),
    .B1(_11120_),
    .C1(_11122_),
    .D1(_10633_),
    .Y(_11129_));
 sky130_fd_sc_hd__o21ai_2 _21296_ (.A1(_11124_),
    .A2(_11126_),
    .B1(net311),
    .Y(_11130_));
 sky130_fd_sc_hd__nand3_1 _21297_ (.A(_11129_),
    .B(net311),
    .C(_11128_),
    .Y(_11131_));
 sky130_fd_sc_hd__o211a_1 _21298_ (.A1(_11100_),
    .A2(net332),
    .B1(_12703_),
    .C1(_11113_),
    .X(_11132_));
 sky130_fd_sc_hd__a211o_1 _21299_ (.A1(_11114_),
    .A2(_11117_),
    .B1(net329),
    .C1(net327),
    .X(_11133_));
 sky130_fd_sc_hd__o22ai_4 _21300_ (.A1(net311),
    .A2(_11119_),
    .B1(_11127_),
    .B2(_11130_),
    .Y(_11134_));
 sky130_fd_sc_hd__a22oi_2 _21301_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_11131_),
    .B2(_11133_),
    .Y(_11135_));
 sky130_fd_sc_hd__o21ai_4 _21302_ (.A1(_06914_),
    .A2(_06916_),
    .B1(_11134_),
    .Y(_11136_));
 sky130_fd_sc_hd__a31oi_1 _21303_ (.A1(_11129_),
    .A2(net311),
    .A3(_11128_),
    .B1(net225),
    .Y(_11137_));
 sky130_fd_sc_hd__a31o_1 _21304_ (.A1(_11129_),
    .A2(net311),
    .A3(_11128_),
    .B1(net225),
    .X(_11138_));
 sky130_fd_sc_hd__o221ai_4 _21305_ (.A1(net311),
    .A2(_11119_),
    .B1(_11127_),
    .B2(_11130_),
    .C1(net227),
    .Y(_11139_));
 sky130_fd_sc_hd__a21oi_1 _21306_ (.A1(_11133_),
    .A2(_11137_),
    .B1(_11135_),
    .Y(_11140_));
 sky130_fd_sc_hd__o21ai_1 _21307_ (.A1(_11132_),
    .A2(_11138_),
    .B1(_11136_),
    .Y(_11141_));
 sky130_fd_sc_hd__o211ai_1 _21308_ (.A1(_09753_),
    .A2(_09759_),
    .B1(_09317_),
    .C1(_09758_),
    .Y(_11142_));
 sky130_fd_sc_hd__nor3_1 _21309_ (.A(_10194_),
    .B(_11142_),
    .C(_10196_),
    .Y(_11143_));
 sky130_fd_sc_hd__nand2_1 _21310_ (.A(_10656_),
    .B(_11143_),
    .Y(_11145_));
 sky130_fd_sc_hd__o211ai_4 _21311_ (.A1(_10661_),
    .A2(_10655_),
    .B1(_10658_),
    .C1(_11145_),
    .Y(_11146_));
 sky130_fd_sc_hd__inv_2 _21312_ (.A(_11146_),
    .Y(_11147_));
 sky130_fd_sc_hd__nand4_4 _21313_ (.A(_11143_),
    .B(_10658_),
    .C(_10656_),
    .D(_09311_),
    .Y(_11148_));
 sky130_fd_sc_hd__inv_2 _21314_ (.A(_11148_),
    .Y(_11149_));
 sky130_fd_sc_hd__nand2_1 _21315_ (.A(_11146_),
    .B(_11148_),
    .Y(_11150_));
 sky130_fd_sc_hd__a21oi_2 _21316_ (.A1(_11146_),
    .A2(_11148_),
    .B1(_11141_),
    .Y(_11151_));
 sky130_fd_sc_hd__o22ai_2 _21317_ (.A1(_00011_),
    .A2(net323),
    .B1(_11140_),
    .B2(_11150_),
    .Y(_11152_));
 sky130_fd_sc_hd__a211o_2 _21318_ (.A1(_11131_),
    .A2(_11133_),
    .B1(_00011_),
    .C1(net323),
    .X(_11153_));
 sky130_fd_sc_hd__inv_2 _21319_ (.A(_11153_),
    .Y(_11154_));
 sky130_fd_sc_hd__nand4_2 _21320_ (.A(_11136_),
    .B(_11139_),
    .C(_11146_),
    .D(_11148_),
    .Y(_11156_));
 sky130_fd_sc_hd__a22o_1 _21321_ (.A1(_11136_),
    .A2(_11139_),
    .B1(_11146_),
    .B2(_11148_),
    .X(_11157_));
 sky130_fd_sc_hd__nand3_2 _21322_ (.A(_11157_),
    .B(net308),
    .C(_11156_),
    .Y(_11158_));
 sky130_fd_sc_hd__o221a_2 _21323_ (.A1(net308),
    .A2(_11134_),
    .B1(_11151_),
    .B2(_11152_),
    .C1(_01973_),
    .X(_11159_));
 sky130_fd_sc_hd__a211o_4 _21324_ (.A1(_11153_),
    .A2(_11158_),
    .B1(net304),
    .C1(_01951_),
    .X(_11160_));
 sky130_fd_sc_hd__a311oi_4 _21325_ (.A1(_11157_),
    .A2(net308),
    .A3(_11156_),
    .B1(net232),
    .C1(_11154_),
    .Y(_11161_));
 sky130_fd_sc_hd__nand3_4 _21326_ (.A(_11158_),
    .B(net234),
    .C(_11153_),
    .Y(_11162_));
 sky130_fd_sc_hd__a2bb2oi_1 _21327_ (.A1_N(_06622_),
    .A2_N(_06624_),
    .B1(_11153_),
    .B2(_11158_),
    .Y(_11163_));
 sky130_fd_sc_hd__o221ai_4 _21328_ (.A1(net308),
    .A2(_11134_),
    .B1(_11151_),
    .B2(_11152_),
    .C1(net232),
    .Y(_11164_));
 sky130_fd_sc_hd__a21oi_1 _21329_ (.A1(net251),
    .A2(_10669_),
    .B1(_10671_),
    .Y(_11165_));
 sky130_fd_sc_hd__o32a_1 _21330_ (.A1(_06305_),
    .A2(_06307_),
    .A3(_10669_),
    .B1(_10671_),
    .B2(_10676_),
    .X(_11167_));
 sky130_fd_sc_hd__a21oi_2 _21331_ (.A1(_10671_),
    .A2(_10675_),
    .B1(_10676_),
    .Y(_11168_));
 sky130_fd_sc_hd__o2bb2ai_4 _21332_ (.A1_N(_11162_),
    .A2_N(_11164_),
    .B1(_11165_),
    .B2(_10674_),
    .Y(_11169_));
 sky130_fd_sc_hd__nand3_4 _21333_ (.A(_11167_),
    .B(_11164_),
    .C(_11162_),
    .Y(_11170_));
 sky130_fd_sc_hd__nand3_4 _21334_ (.A(_11169_),
    .B(_11170_),
    .C(net279),
    .Y(_11171_));
 sky130_fd_sc_hd__a31o_2 _21335_ (.A1(_11169_),
    .A2(_11170_),
    .A3(net279),
    .B1(_11159_),
    .X(_11172_));
 sky130_fd_sc_hd__o21ai_4 _21336_ (.A1(net254),
    .A2(_10689_),
    .B1(_10697_),
    .Y(_11173_));
 sky130_fd_sc_hd__a22oi_1 _21337_ (.A1(net254),
    .A2(_10689_),
    .B1(_10228_),
    .B2(_10219_),
    .Y(_11174_));
 sky130_fd_sc_hd__a22o_1 _21338_ (.A1(net254),
    .A2(_10689_),
    .B1(_10228_),
    .B2(_10219_),
    .X(_11175_));
 sky130_fd_sc_hd__a31oi_2 _21339_ (.A1(_11169_),
    .A2(_11170_),
    .A3(net279),
    .B1(net251),
    .Y(_11176_));
 sky130_fd_sc_hd__a311oi_4 _21340_ (.A1(_11169_),
    .A2(_11170_),
    .A3(net279),
    .B1(net251),
    .C1(_11159_),
    .Y(_11178_));
 sky130_fd_sc_hd__o211ai_4 _21341_ (.A1(_06309_),
    .A2(_06312_),
    .B1(_11160_),
    .C1(_11171_),
    .Y(_11179_));
 sky130_fd_sc_hd__a2bb2oi_4 _21342_ (.A1_N(_06305_),
    .A2_N(_06307_),
    .B1(_11160_),
    .B2(_11171_),
    .Y(_11180_));
 sky130_fd_sc_hd__a22o_1 _21343_ (.A1(_06306_),
    .A2(_06308_),
    .B1(_11160_),
    .B2(_11171_),
    .X(_11181_));
 sky130_fd_sc_hd__o2111ai_1 _21344_ (.A1(_10689_),
    .A2(net254),
    .B1(_11179_),
    .C1(_11175_),
    .D1(_11181_),
    .Y(_11182_));
 sky130_fd_sc_hd__o22ai_1 _21345_ (.A1(_10690_),
    .A2(_11174_),
    .B1(_11178_),
    .B2(_11180_),
    .Y(_11183_));
 sky130_fd_sc_hd__o2111ai_2 _21346_ (.A1(net253),
    .A2(_10688_),
    .B1(_11173_),
    .C1(_11179_),
    .D1(_11181_),
    .Y(_11184_));
 sky130_fd_sc_hd__o2bb2ai_1 _21347_ (.A1_N(_10693_),
    .A2_N(_11173_),
    .B1(_11178_),
    .B2(_11180_),
    .Y(_11185_));
 sky130_fd_sc_hd__nand3_2 _21348_ (.A(_11182_),
    .B(_11183_),
    .C(net277),
    .Y(_11186_));
 sky130_fd_sc_hd__a21oi_1 _21349_ (.A1(_11160_),
    .A2(_11171_),
    .B1(net277),
    .Y(_11187_));
 sky130_fd_sc_hd__nand3_1 _21350_ (.A(_11184_),
    .B(_11185_),
    .C(net277),
    .Y(_11189_));
 sky130_fd_sc_hd__a31o_1 _21351_ (.A1(_11184_),
    .A2(_11185_),
    .A3(net277),
    .B1(_11187_),
    .X(_11190_));
 sky130_fd_sc_hd__o21ai_4 _21352_ (.A1(net277),
    .A2(_11172_),
    .B1(_11186_),
    .Y(_11191_));
 sky130_fd_sc_hd__o21a_1 _21353_ (.A1(_05228_),
    .A2(_05230_),
    .B1(_11191_),
    .X(_11192_));
 sky130_fd_sc_hd__a311o_1 _21354_ (.A1(_11184_),
    .A2(_11185_),
    .A3(net277),
    .B1(_11187_),
    .C1(net272),
    .X(_11193_));
 sky130_fd_sc_hd__nand3b_4 _21355_ (.A_N(_11187_),
    .B(_11189_),
    .C(net254),
    .Y(_11194_));
 sky130_fd_sc_hd__o211ai_4 _21356_ (.A1(_11172_),
    .A2(net276),
    .B1(net253),
    .C1(_11186_),
    .Y(_11195_));
 sky130_fd_sc_hd__nand2_1 _21357_ (.A(_11194_),
    .B(_11195_),
    .Y(_11196_));
 sky130_fd_sc_hd__o2bb2ai_2 _21358_ (.A1_N(_10710_),
    .A2_N(_10712_),
    .B1(net262),
    .B2(_10705_),
    .Y(_11197_));
 sky130_fd_sc_hd__o211ai_4 _21359_ (.A1(_10239_),
    .A2(_10711_),
    .B1(_10719_),
    .C1(_10710_),
    .Y(_11198_));
 sky130_fd_sc_hd__o2111ai_4 _21360_ (.A1(_10705_),
    .A2(net262),
    .B1(_11195_),
    .C1(_11194_),
    .D1(_11198_),
    .Y(_11200_));
 sky130_fd_sc_hd__a22o_1 _21361_ (.A1(_11194_),
    .A2(_11195_),
    .B1(_11198_),
    .B2(_10715_),
    .X(_11201_));
 sky130_fd_sc_hd__o211ai_1 _21362_ (.A1(_05231_),
    .A2(_05232_),
    .B1(_11200_),
    .C1(_11201_),
    .Y(_11202_));
 sky130_fd_sc_hd__o211a_1 _21363_ (.A1(_11172_),
    .A2(net276),
    .B1(_05234_),
    .C1(_11186_),
    .X(_11203_));
 sky130_fd_sc_hd__o211ai_2 _21364_ (.A1(_10705_),
    .A2(net262),
    .B1(_11198_),
    .C1(_11196_),
    .Y(_11204_));
 sky130_fd_sc_hd__o2111ai_4 _21365_ (.A1(net261),
    .A2(_10704_),
    .B1(_11194_),
    .C1(_11195_),
    .D1(_11197_),
    .Y(_11205_));
 sky130_fd_sc_hd__o211a_1 _21366_ (.A1(_05231_),
    .A2(_05232_),
    .B1(_11204_),
    .C1(_11205_),
    .X(_11206_));
 sky130_fd_sc_hd__o211ai_2 _21367_ (.A1(_05231_),
    .A2(_05232_),
    .B1(_11204_),
    .C1(_11205_),
    .Y(_11207_));
 sky130_fd_sc_hd__a31o_2 _21368_ (.A1(_11204_),
    .A2(_11205_),
    .A3(net272),
    .B1(_11203_),
    .X(_11208_));
 sky130_fd_sc_hd__a31o_1 _21369_ (.A1(_11201_),
    .A2(net273),
    .A3(_11200_),
    .B1(_11192_),
    .X(_11209_));
 sky130_fd_sc_hd__and3_1 _21370_ (.A(net261),
    .B(_11193_),
    .C(_11202_),
    .X(_11211_));
 sky130_fd_sc_hd__a311o_2 _21371_ (.A1(_11201_),
    .A2(net273),
    .A3(_11200_),
    .B1(net262),
    .C1(_11192_),
    .X(_11212_));
 sky130_fd_sc_hd__o221ai_4 _21372_ (.A1(_05765_),
    .A2(net289),
    .B1(_11191_),
    .B2(net273),
    .C1(_11207_),
    .Y(_11213_));
 sky130_fd_sc_hd__nand2_1 _21373_ (.A(_11212_),
    .B(_11213_),
    .Y(_11214_));
 sky130_fd_sc_hd__nand4_2 _21374_ (.A(_09375_),
    .B(_09377_),
    .C(_09836_),
    .D(_09838_),
    .Y(_11215_));
 sky130_fd_sc_hd__a21oi_1 _21375_ (.A1(net294),
    .A2(_10252_),
    .B1(_11215_),
    .Y(_11216_));
 sky130_fd_sc_hd__nor3_2 _21376_ (.A(_11215_),
    .B(_10260_),
    .C(_10258_),
    .Y(_11217_));
 sky130_fd_sc_hd__o211ai_2 _21377_ (.A1(net294),
    .A2(_10252_),
    .B1(_11216_),
    .C1(_10734_),
    .Y(_11218_));
 sky130_fd_sc_hd__o2111ai_2 _21378_ (.A1(net294),
    .A2(_10252_),
    .B1(_11216_),
    .C1(_10734_),
    .D1(_09385_),
    .Y(_11219_));
 sky130_fd_sc_hd__o221ai_4 _21379_ (.A1(_10729_),
    .A2(net292),
    .B1(_11217_),
    .B2(_10742_),
    .C1(_11219_),
    .Y(_11220_));
 sky130_fd_sc_hd__o211ai_4 _21380_ (.A1(_10740_),
    .A2(_10733_),
    .B1(_10735_),
    .C1(_11218_),
    .Y(_11222_));
 sky130_fd_sc_hd__nand4_4 _21381_ (.A(_11217_),
    .B(_10735_),
    .C(_10734_),
    .D(_09385_),
    .Y(_11223_));
 sky130_fd_sc_hd__o21a_2 _21382_ (.A1(net267),
    .A2(_10730_),
    .B1(_11220_),
    .X(_11224_));
 sky130_fd_sc_hd__inv_2 _21383_ (.A(_11224_),
    .Y(_11225_));
 sky130_fd_sc_hd__o211ai_4 _21384_ (.A1(net267),
    .A2(_10730_),
    .B1(_11214_),
    .C1(_11220_),
    .Y(_11226_));
 sky130_fd_sc_hd__o31a_1 _21385_ (.A1(net261),
    .A2(_11203_),
    .A3(_11206_),
    .B1(_11223_),
    .X(_11227_));
 sky130_fd_sc_hd__o211ai_2 _21386_ (.A1(_11208_),
    .A2(net261),
    .B1(_11223_),
    .C1(_11222_),
    .Y(_11228_));
 sky130_fd_sc_hd__o2111ai_4 _21387_ (.A1(net261),
    .A2(_11208_),
    .B1(_11212_),
    .C1(_11222_),
    .D1(_11223_),
    .Y(_11229_));
 sky130_fd_sc_hd__nand3_2 _21388_ (.A(_11226_),
    .B(_11229_),
    .C(net246),
    .Y(_11230_));
 sky130_fd_sc_hd__and3_4 _21389_ (.A(_05486_),
    .B(_11193_),
    .C(_11202_),
    .X(_11231_));
 sky130_fd_sc_hd__a311o_2 _21390_ (.A1(_11201_),
    .A2(net273),
    .A3(_11200_),
    .B1(net246),
    .C1(_11192_),
    .X(_11233_));
 sky130_fd_sc_hd__a31oi_4 _21391_ (.A1(_11226_),
    .A2(_11229_),
    .A3(net246),
    .B1(_11231_),
    .Y(_11234_));
 sky130_fd_sc_hd__a21oi_4 _21392_ (.A1(_11230_),
    .A2(_11233_),
    .B1(net242),
    .Y(_11235_));
 sky130_fd_sc_hd__or3_1 _21393_ (.A(net266),
    .B(_05751_),
    .C(_11234_),
    .X(_11236_));
 sky130_fd_sc_hd__a31o_2 _21394_ (.A1(_11226_),
    .A2(_11229_),
    .A3(net246),
    .B1(net291),
    .X(_11237_));
 sky130_fd_sc_hd__a311oi_4 _21395_ (.A1(_11226_),
    .A2(_11229_),
    .A3(net246),
    .B1(_11231_),
    .C1(net292),
    .Y(_11238_));
 sky130_fd_sc_hd__a31o_1 _21396_ (.A1(_05482_),
    .A2(_05484_),
    .A3(_11208_),
    .B1(_11237_),
    .X(_11239_));
 sky130_fd_sc_hd__a22oi_4 _21397_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_11230_),
    .B2(_11233_),
    .Y(_11240_));
 sky130_fd_sc_hd__a21o_1 _21398_ (.A1(_11230_),
    .A2(_11233_),
    .B1(net267),
    .X(_11241_));
 sky130_fd_sc_hd__o32a_2 _21399_ (.A1(net318),
    .A2(_05244_),
    .A3(_10745_),
    .B1(_10748_),
    .B2(_10752_),
    .X(_11242_));
 sky130_fd_sc_hd__a21oi_2 _21400_ (.A1(_10751_),
    .A2(_10748_),
    .B1(_10752_),
    .Y(_11244_));
 sky130_fd_sc_hd__o21a_1 _21401_ (.A1(_11238_),
    .A2(_11240_),
    .B1(_11244_),
    .X(_11245_));
 sky130_fd_sc_hd__o21ai_4 _21402_ (.A1(_11238_),
    .A2(_11240_),
    .B1(_11244_),
    .Y(_11246_));
 sky130_fd_sc_hd__o21ai_1 _21403_ (.A1(net267),
    .A2(_11234_),
    .B1(_11242_),
    .Y(_11247_));
 sky130_fd_sc_hd__o211ai_4 _21404_ (.A1(_11231_),
    .A2(_11237_),
    .B1(_11242_),
    .C1(_11241_),
    .Y(_11248_));
 sky130_fd_sc_hd__o22ai_2 _21405_ (.A1(net266),
    .A2(_05751_),
    .B1(_11238_),
    .B2(_11247_),
    .Y(_11249_));
 sky130_fd_sc_hd__o211ai_2 _21406_ (.A1(_11238_),
    .A2(_11247_),
    .B1(net242),
    .C1(_11246_),
    .Y(_11250_));
 sky130_fd_sc_hd__a31oi_4 _21407_ (.A1(_11246_),
    .A2(_11248_),
    .A3(net242),
    .B1(_11235_),
    .Y(_11251_));
 sky130_fd_sc_hd__o22ai_4 _21408_ (.A1(net242),
    .A2(_11234_),
    .B1(_11245_),
    .B2(_11249_),
    .Y(_11252_));
 sky130_fd_sc_hd__a311o_1 _21409_ (.A1(_11246_),
    .A2(_11248_),
    .A3(net242),
    .B1(net240),
    .C1(_11235_),
    .X(_11253_));
 sky130_fd_sc_hd__o311a_1 _21410_ (.A1(_10293_),
    .A2(_10301_),
    .A3(_10304_),
    .B1(_10765_),
    .C1(_10291_),
    .X(_11255_));
 sky130_fd_sc_hd__a21oi_1 _21411_ (.A1(_10291_),
    .A2(_10315_),
    .B1(_10766_),
    .Y(_11256_));
 sky130_fd_sc_hd__a21o_1 _21412_ (.A1(_10769_),
    .A2(_10767_),
    .B1(_10764_),
    .X(_11257_));
 sky130_fd_sc_hd__a31o_1 _21413_ (.A1(_11246_),
    .A2(_11248_),
    .A3(net242),
    .B1(net294),
    .X(_11258_));
 sky130_fd_sc_hd__a311oi_4 _21414_ (.A1(_11246_),
    .A2(_11248_),
    .A3(net242),
    .B1(_11235_),
    .C1(net294),
    .Y(_11259_));
 sky130_fd_sc_hd__nand3_2 _21415_ (.A(_11250_),
    .B(net295),
    .C(_11236_),
    .Y(_11260_));
 sky130_fd_sc_hd__a2bb2oi_2 _21416_ (.A1_N(net318),
    .A2_N(_05244_),
    .B1(_11236_),
    .B2(_11250_),
    .Y(_11261_));
 sky130_fd_sc_hd__o21ai_4 _21417_ (.A1(net318),
    .A2(net316),
    .B1(_11252_),
    .Y(_11262_));
 sky130_fd_sc_hd__o221ai_2 _21418_ (.A1(_10766_),
    .A2(_11255_),
    .B1(_11235_),
    .B2(_11258_),
    .C1(_11262_),
    .Y(_11263_));
 sky130_fd_sc_hd__o22ai_1 _21419_ (.A1(_10764_),
    .A2(_11256_),
    .B1(_11259_),
    .B2(_11261_),
    .Y(_11264_));
 sky130_fd_sc_hd__o211ai_2 _21420_ (.A1(net259),
    .A2(_05992_),
    .B1(_11263_),
    .C1(_11264_),
    .Y(_11266_));
 sky130_fd_sc_hd__or3_1 _21421_ (.A(_05990_),
    .B(_05992_),
    .C(_11251_),
    .X(_11267_));
 sky130_fd_sc_hd__o21ai_1 _21422_ (.A1(net295),
    .A2(_11251_),
    .B1(_11257_),
    .Y(_11268_));
 sky130_fd_sc_hd__o22ai_2 _21423_ (.A1(_10766_),
    .A2(_11255_),
    .B1(_11259_),
    .B2(_11261_),
    .Y(_11269_));
 sky130_fd_sc_hd__o221ai_4 _21424_ (.A1(net259),
    .A2(_05992_),
    .B1(_11259_),
    .B2(_11268_),
    .C1(_11269_),
    .Y(_11270_));
 sky130_fd_sc_hd__o21ai_1 _21425_ (.A1(net240),
    .A2(_11251_),
    .B1(_11270_),
    .Y(_11271_));
 sky130_fd_sc_hd__o31a_1 _21426_ (.A1(_05990_),
    .A2(_05992_),
    .A3(_11251_),
    .B1(_11270_),
    .X(_11272_));
 sky130_fd_sc_hd__o211ai_4 _21427_ (.A1(net341),
    .A2(_04184_),
    .B1(_11253_),
    .C1(_11266_),
    .Y(_11273_));
 sky130_fd_sc_hd__o311a_1 _21428_ (.A1(_05990_),
    .A2(_05992_),
    .A3(_11251_),
    .B1(net299),
    .C1(_11270_),
    .X(_11274_));
 sky130_fd_sc_hd__o211ai_2 _21429_ (.A1(net240),
    .A2(_11251_),
    .B1(net299),
    .C1(_11270_),
    .Y(_11275_));
 sky130_fd_sc_hd__a21oi_1 _21430_ (.A1(_10790_),
    .A2(_10793_),
    .B1(_10777_),
    .Y(_11277_));
 sky130_fd_sc_hd__a31oi_2 _21431_ (.A1(_10781_),
    .A2(_10790_),
    .A3(_10793_),
    .B1(_10777_),
    .Y(_11278_));
 sky130_fd_sc_hd__o2bb2ai_1 _21432_ (.A1_N(_02148_),
    .A2_N(_10776_),
    .B1(_10789_),
    .B2(_10796_),
    .Y(_11279_));
 sky130_fd_sc_hd__o2bb2ai_1 _21433_ (.A1_N(_11273_),
    .A2_N(_11275_),
    .B1(_11277_),
    .B2(_10780_),
    .Y(_11280_));
 sky130_fd_sc_hd__nand3_1 _21434_ (.A(_11273_),
    .B(_11275_),
    .C(_11279_),
    .Y(_11281_));
 sky130_fd_sc_hd__o311a_1 _21435_ (.A1(_05990_),
    .A2(_11252_),
    .A3(_05992_),
    .B1(_06294_),
    .C1(_11266_),
    .X(_11282_));
 sky130_fd_sc_hd__a22o_1 _21436_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_11267_),
    .B2(_11270_),
    .X(_11283_));
 sky130_fd_sc_hd__nand3_1 _21437_ (.A(_11280_),
    .B(_11281_),
    .C(net213),
    .Y(_11284_));
 sky130_fd_sc_hd__a31o_2 _21438_ (.A1(_11280_),
    .A2(_11281_),
    .A3(net213),
    .B1(_11282_),
    .X(_11285_));
 sky130_fd_sc_hd__o31a_1 _21439_ (.A1(_06291_),
    .A2(_06292_),
    .A3(_11272_),
    .B1(_11284_),
    .X(_11286_));
 sky130_fd_sc_hd__a21oi_1 _21440_ (.A1(_11283_),
    .A2(_11284_),
    .B1(_02137_),
    .Y(_11288_));
 sky130_fd_sc_hd__a22o_1 _21441_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_11283_),
    .B2(_11284_),
    .X(_11289_));
 sky130_fd_sc_hd__and3_1 _21442_ (.A(_11284_),
    .B(_02137_),
    .C(_11283_),
    .X(_11290_));
 sky130_fd_sc_hd__a311o_1 _21443_ (.A1(_11280_),
    .A2(_11281_),
    .A3(net213),
    .B1(_11282_),
    .C1(_02148_),
    .X(_11291_));
 sky130_fd_sc_hd__nand4_1 _21444_ (.A(_09449_),
    .B(_09451_),
    .C(_09904_),
    .D(_09906_),
    .Y(_11292_));
 sky130_fd_sc_hd__nor3_1 _21445_ (.A(_10340_),
    .B(_11292_),
    .C(_10342_),
    .Y(_11293_));
 sky130_fd_sc_hd__nand2_1 _21446_ (.A(_10809_),
    .B(_11293_),
    .Y(_11294_));
 sky130_fd_sc_hd__o211ai_4 _21447_ (.A1(_10813_),
    .A2(_10808_),
    .B1(_10811_),
    .C1(_11294_),
    .Y(_11295_));
 sky130_fd_sc_hd__nor4_1 _21448_ (.A(_09454_),
    .B(_11292_),
    .C(_10342_),
    .D(_10340_),
    .Y(_11296_));
 sky130_fd_sc_hd__o211ai_2 _21449_ (.A1(_00240_),
    .A2(_10803_),
    .B1(_11293_),
    .C1(_09453_),
    .Y(_11297_));
 sky130_fd_sc_hd__nand3_4 _21450_ (.A(_10809_),
    .B(_10811_),
    .C(_11296_),
    .Y(_11299_));
 sky130_fd_sc_hd__o21ai_4 _21451_ (.A1(_10808_),
    .A2(_11297_),
    .B1(_11295_),
    .Y(_11300_));
 sky130_fd_sc_hd__o21ai_4 _21452_ (.A1(_11288_),
    .A2(_11290_),
    .B1(_11300_),
    .Y(_11301_));
 sky130_fd_sc_hd__o211ai_2 _21453_ (.A1(_02148_),
    .A2(_11285_),
    .B1(_11295_),
    .C1(_11299_),
    .Y(_11302_));
 sky130_fd_sc_hd__nand4_4 _21454_ (.A(_11289_),
    .B(_11291_),
    .C(_11295_),
    .D(_11299_),
    .Y(_11303_));
 sky130_fd_sc_hd__nand3_2 _21455_ (.A(_11301_),
    .B(_11303_),
    .C(net211),
    .Y(_11304_));
 sky130_fd_sc_hd__and3_4 _21456_ (.A(_11285_),
    .B(_06611_),
    .C(_06609_),
    .X(_11305_));
 sky130_fd_sc_hd__or3_2 _21457_ (.A(_06608_),
    .B(net237),
    .C(_11286_),
    .X(_11306_));
 sky130_fd_sc_hd__a31oi_4 _21458_ (.A1(_11301_),
    .A2(_11303_),
    .A3(net211),
    .B1(_11305_),
    .Y(_11307_));
 sky130_fd_sc_hd__a21oi_2 _21459_ (.A1(_11304_),
    .A2(_11306_),
    .B1(net208),
    .Y(_11308_));
 sky130_fd_sc_hd__or3_2 _21460_ (.A(net230),
    .B(_06901_),
    .C(_11307_),
    .X(_11310_));
 sky130_fd_sc_hd__a31o_1 _21461_ (.A1(_11301_),
    .A2(_11303_),
    .A3(net211),
    .B1(_00251_),
    .X(_11311_));
 sky130_fd_sc_hd__a311oi_4 _21462_ (.A1(_11301_),
    .A2(_11303_),
    .A3(net211),
    .B1(_11305_),
    .C1(_00251_),
    .Y(_11312_));
 sky130_fd_sc_hd__a311o_1 _21463_ (.A1(_11301_),
    .A2(_11303_),
    .A3(net211),
    .B1(_11305_),
    .C1(_00251_),
    .X(_11313_));
 sky130_fd_sc_hd__a22oi_4 _21464_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_11304_),
    .B2(_11306_),
    .Y(_11314_));
 sky130_fd_sc_hd__a22o_1 _21465_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_11304_),
    .B2(_11306_),
    .X(_11315_));
 sky130_fd_sc_hd__a21o_2 _21466_ (.A1(_10823_),
    .A2(_10821_),
    .B1(_10824_),
    .X(_11316_));
 sky130_fd_sc_hd__o31a_1 _21467_ (.A1(_10356_),
    .A2(_10820_),
    .A3(_10822_),
    .B1(_10825_),
    .X(_11317_));
 sky130_fd_sc_hd__o21a_1 _21468_ (.A1(_11312_),
    .A2(_11314_),
    .B1(_11317_),
    .X(_11318_));
 sky130_fd_sc_hd__o21ai_4 _21469_ (.A1(_11312_),
    .A2(_11314_),
    .B1(_11317_),
    .Y(_11319_));
 sky130_fd_sc_hd__o21ai_2 _21470_ (.A1(_00240_),
    .A2(_11307_),
    .B1(_11316_),
    .Y(_11321_));
 sky130_fd_sc_hd__o211ai_4 _21471_ (.A1(_11305_),
    .A2(_11311_),
    .B1(_11316_),
    .C1(_11315_),
    .Y(_11322_));
 sky130_fd_sc_hd__o22ai_2 _21472_ (.A1(net230),
    .A2(_06901_),
    .B1(_11312_),
    .B2(_11321_),
    .Y(_11323_));
 sky130_fd_sc_hd__o211ai_4 _21473_ (.A1(_11312_),
    .A2(_11321_),
    .B1(net208),
    .C1(_11319_),
    .Y(_11324_));
 sky130_fd_sc_hd__o22ai_4 _21474_ (.A1(net208),
    .A2(_11307_),
    .B1(_11318_),
    .B2(_11323_),
    .Y(_11325_));
 sky130_fd_sc_hd__a311o_2 _21475_ (.A1(_11319_),
    .A2(_11322_),
    .A3(net208),
    .B1(net185),
    .C1(_11308_),
    .X(_11326_));
 sky130_fd_sc_hd__o311a_1 _21476_ (.A1(net365),
    .A2(net362),
    .A3(_10365_),
    .B1(_10374_),
    .C1(_10840_),
    .X(_11327_));
 sky130_fd_sc_hd__o32a_1 _21477_ (.A1(_11309_),
    .A2(_10830_),
    .A3(_10834_),
    .B1(_10367_),
    .B2(_10373_),
    .X(_11328_));
 sky130_fd_sc_hd__a21o_1 _21478_ (.A1(_10842_),
    .A2(_10843_),
    .B1(_10839_),
    .X(_11329_));
 sky130_fd_sc_hd__a21oi_1 _21479_ (.A1(_10842_),
    .A2(_10843_),
    .B1(_10839_),
    .Y(_11330_));
 sky130_fd_sc_hd__a31oi_1 _21480_ (.A1(_11319_),
    .A2(_11322_),
    .A3(net208),
    .B1(net326),
    .Y(_11332_));
 sky130_fd_sc_hd__a311oi_4 _21481_ (.A1(_11319_),
    .A2(_11322_),
    .A3(net208),
    .B1(_11308_),
    .C1(net326),
    .Y(_11333_));
 sky130_fd_sc_hd__o221ai_4 _21482_ (.A1(_12867_),
    .A2(_12877_),
    .B1(net208),
    .B2(_11307_),
    .C1(_11324_),
    .Y(_11334_));
 sky130_fd_sc_hd__a2bb2oi_2 _21483_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_11310_),
    .B2(_11324_),
    .Y(_11335_));
 sky130_fd_sc_hd__o21ai_2 _21484_ (.A1(net361),
    .A2(net345),
    .B1(_11325_),
    .Y(_11336_));
 sky130_fd_sc_hd__o211ai_2 _21485_ (.A1(_10841_),
    .A2(_11327_),
    .B1(_11334_),
    .C1(_11336_),
    .Y(_11337_));
 sky130_fd_sc_hd__o22ai_2 _21486_ (.A1(_10839_),
    .A2(_11328_),
    .B1(_11333_),
    .B2(_11335_),
    .Y(_11338_));
 sky130_fd_sc_hd__o211ai_4 _21487_ (.A1(_07227_),
    .A2(_07229_),
    .B1(_11337_),
    .C1(_11338_),
    .Y(_11339_));
 sky130_fd_sc_hd__a211o_2 _21488_ (.A1(_11310_),
    .A2(_11324_),
    .B1(_07227_),
    .C1(net203),
    .X(_11340_));
 sky130_fd_sc_hd__o211ai_2 _21489_ (.A1(_10839_),
    .A2(_11328_),
    .B1(_11334_),
    .C1(_11336_),
    .Y(_11341_));
 sky130_fd_sc_hd__o22ai_2 _21490_ (.A1(_10841_),
    .A2(_11327_),
    .B1(_11333_),
    .B2(_11335_),
    .Y(_11343_));
 sky130_fd_sc_hd__o211ai_4 _21491_ (.A1(_07227_),
    .A2(net203),
    .B1(_11341_),
    .C1(_11343_),
    .Y(_11344_));
 sky130_fd_sc_hd__o21ai_4 _21492_ (.A1(net185),
    .A2(_11325_),
    .B1(_11339_),
    .Y(_11345_));
 sky130_fd_sc_hd__a2bb2oi_1 _21493_ (.A1_N(_11210_),
    .A2_N(_11232_),
    .B1(_11340_),
    .B2(_11344_),
    .Y(_11346_));
 sky130_fd_sc_hd__o211ai_4 _21494_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_11326_),
    .C1(_11339_),
    .Y(_11347_));
 sky130_fd_sc_hd__o211ai_4 _21495_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_11340_),
    .C1(_11344_),
    .Y(_11348_));
 sky130_fd_sc_hd__o211a_1 _21496_ (.A1(_10383_),
    .A2(_10384_),
    .B1(_10387_),
    .C1(_10851_),
    .X(_11349_));
 sky130_fd_sc_hd__nand2_2 _21497_ (.A(_10851_),
    .B(_10859_),
    .Y(_11350_));
 sky130_fd_sc_hd__a21oi_2 _21498_ (.A1(_11347_),
    .A2(_11348_),
    .B1(_11350_),
    .Y(_11351_));
 sky130_fd_sc_hd__o2bb2ai_1 _21499_ (.A1_N(_11347_),
    .A2_N(_11348_),
    .B1(_11349_),
    .B2(_10853_),
    .Y(_11352_));
 sky130_fd_sc_hd__nand3_1 _21500_ (.A(_11347_),
    .B(_11348_),
    .C(_11350_),
    .Y(_11354_));
 sky130_fd_sc_hd__a31o_1 _21501_ (.A1(_11347_),
    .A2(_11348_),
    .A3(_11350_),
    .B1(_07550_),
    .X(_11355_));
 sky130_fd_sc_hd__nand3_2 _21502_ (.A(_11352_),
    .B(_11354_),
    .C(net163),
    .Y(_11356_));
 sky130_fd_sc_hd__a211o_1 _21503_ (.A1(_11340_),
    .A2(_11344_),
    .B1(_07544_),
    .C1(net184),
    .X(_11357_));
 sky130_fd_sc_hd__o32a_2 _21504_ (.A1(_07544_),
    .A2(net184),
    .A3(_11345_),
    .B1(_11351_),
    .B2(_11355_),
    .X(_11358_));
 sky130_fd_sc_hd__o22ai_4 _21505_ (.A1(net163),
    .A2(_11345_),
    .B1(_11351_),
    .B2(_11355_),
    .Y(_11359_));
 sky130_fd_sc_hd__and3_1 _21506_ (.A(_07913_),
    .B(_07915_),
    .C(_11359_),
    .X(_11360_));
 sky130_fd_sc_hd__or3_2 _21507_ (.A(_07912_),
    .B(_07914_),
    .C(_11358_),
    .X(_11361_));
 sky130_fd_sc_hd__o31a_2 _21508_ (.A1(_10864_),
    .A2(_08918_),
    .A3(_10862_),
    .B1(_10868_),
    .X(_11362_));
 sky130_fd_sc_hd__a21o_2 _21509_ (.A1(_10868_),
    .A2(_10870_),
    .B1(_10872_),
    .X(_11363_));
 sky130_fd_sc_hd__a22oi_4 _21510_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_11356_),
    .B2(_11357_),
    .Y(_11365_));
 sky130_fd_sc_hd__o21ai_2 _21511_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_11359_),
    .Y(_11366_));
 sky130_fd_sc_hd__o221a_1 _21512_ (.A1(net163),
    .A2(_11345_),
    .B1(_11351_),
    .B2(_11355_),
    .C1(_10015_),
    .X(_11367_));
 sky130_fd_sc_hd__o221ai_4 _21513_ (.A1(net365),
    .A2(net362),
    .B1(net163),
    .B2(_11345_),
    .C1(_11356_),
    .Y(_11368_));
 sky130_fd_sc_hd__a21oi_2 _21514_ (.A1(_11366_),
    .A2(_11368_),
    .B1(_11363_),
    .Y(_11369_));
 sky130_fd_sc_hd__o21bai_4 _21515_ (.A1(_11365_),
    .A2(_11367_),
    .B1_N(_11363_),
    .Y(_11370_));
 sky130_fd_sc_hd__o21ai_4 _21516_ (.A1(_10872_),
    .A2(_11362_),
    .B1(_11368_),
    .Y(_11371_));
 sky130_fd_sc_hd__o221ai_4 _21517_ (.A1(_10025_),
    .A2(_11359_),
    .B1(_11362_),
    .B2(_10872_),
    .C1(_11366_),
    .Y(_11372_));
 sky130_fd_sc_hd__o22ai_4 _21518_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_11365_),
    .B2(_11371_),
    .Y(_11373_));
 sky130_fd_sc_hd__o211ai_4 _21519_ (.A1(_11365_),
    .A2(_11371_),
    .B1(net160),
    .C1(_11370_),
    .Y(_11374_));
 sky130_fd_sc_hd__o22ai_2 _21520_ (.A1(net160),
    .A2(_11358_),
    .B1(_11369_),
    .B2(_11373_),
    .Y(_11376_));
 sky130_fd_sc_hd__and3_2 _21521_ (.A(_08297_),
    .B(_08299_),
    .C(_11376_),
    .X(_11377_));
 sky130_fd_sc_hd__a211o_1 _21522_ (.A1(_11361_),
    .A2(_11374_),
    .B1(net180),
    .C1(_08298_),
    .X(_11378_));
 sky130_fd_sc_hd__a21oi_2 _21523_ (.A1(_07899_),
    .A2(_10877_),
    .B1(_10880_),
    .Y(_11379_));
 sky130_fd_sc_hd__o32a_1 _21524_ (.A1(_07800_),
    .A2(_07822_),
    .A3(_10877_),
    .B1(_10880_),
    .B2(_10884_),
    .X(_11380_));
 sky130_fd_sc_hd__a311oi_4 _21525_ (.A1(_11370_),
    .A2(_11372_),
    .A3(net160),
    .B1(_11360_),
    .C1(_08918_),
    .Y(_11381_));
 sky130_fd_sc_hd__o221ai_4 _21526_ (.A1(net160),
    .A2(_11358_),
    .B1(_11369_),
    .B2(_11373_),
    .C1(_08907_),
    .Y(_11382_));
 sky130_fd_sc_hd__a2bb2oi_4 _21527_ (.A1_N(_08819_),
    .A2_N(_08841_),
    .B1(_11361_),
    .B2(_11374_),
    .Y(_11383_));
 sky130_fd_sc_hd__o21ai_2 _21528_ (.A1(_08819_),
    .A2(_08841_),
    .B1(_11376_),
    .Y(_11384_));
 sky130_fd_sc_hd__o22ai_1 _21529_ (.A1(_10884_),
    .A2(_10890_),
    .B1(_11381_),
    .B2(_11383_),
    .Y(_11385_));
 sky130_fd_sc_hd__o211ai_1 _21530_ (.A1(_10881_),
    .A2(_11379_),
    .B1(_11382_),
    .C1(_11384_),
    .Y(_11387_));
 sky130_fd_sc_hd__o211ai_4 _21531_ (.A1(_10884_),
    .A2(_10890_),
    .B1(_11382_),
    .C1(_11384_),
    .Y(_11388_));
 sky130_fd_sc_hd__o22ai_4 _21532_ (.A1(_10881_),
    .A2(_11379_),
    .B1(_11381_),
    .B2(_11383_),
    .Y(_11389_));
 sky130_fd_sc_hd__a22oi_2 _21533_ (.A1(_08297_),
    .A2(_08299_),
    .B1(_11385_),
    .B2(_11387_),
    .Y(_11390_));
 sky130_fd_sc_hd__o211ai_2 _21534_ (.A1(net180),
    .A2(_08298_),
    .B1(_11388_),
    .C1(_11389_),
    .Y(_11391_));
 sky130_fd_sc_hd__a31o_1 _21535_ (.A1(_11389_),
    .A2(_08300_),
    .A3(_11388_),
    .B1(_11377_),
    .X(_11392_));
 sky130_fd_sc_hd__and3_1 _21536_ (.A(_08710_),
    .B(_08713_),
    .C(_11392_),
    .X(_11393_));
 sky130_fd_sc_hd__a22o_1 _21537_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_11378_),
    .B2(_11391_),
    .X(_11394_));
 sky130_fd_sc_hd__o311a_1 _21538_ (.A1(_09996_),
    .A2(_10431_),
    .A3(_10434_),
    .B1(_10899_),
    .C1(_10430_),
    .X(_11395_));
 sky130_fd_sc_hd__a21o_1 _21539_ (.A1(_10484_),
    .A2(_10896_),
    .B1(_10898_),
    .X(_11396_));
 sky130_fd_sc_hd__a21oi_1 _21540_ (.A1(_10484_),
    .A2(_10896_),
    .B1(_10898_),
    .Y(_11398_));
 sky130_fd_sc_hd__a311oi_4 _21541_ (.A1(_11388_),
    .A2(_11389_),
    .A3(_08300_),
    .B1(_11377_),
    .C1(_07899_),
    .Y(_11399_));
 sky130_fd_sc_hd__o211ai_1 _21542_ (.A1(net368),
    .A2(_07866_),
    .B1(_11378_),
    .C1(_11391_),
    .Y(_11400_));
 sky130_fd_sc_hd__a21oi_2 _21543_ (.A1(_11378_),
    .A2(_11391_),
    .B1(_07888_),
    .Y(_11401_));
 sky130_fd_sc_hd__o22ai_2 _21544_ (.A1(_07800_),
    .A2(_07822_),
    .B1(_11377_),
    .B2(_11390_),
    .Y(_11402_));
 sky130_fd_sc_hd__o31a_1 _21545_ (.A1(_07899_),
    .A2(_11377_),
    .A3(_11390_),
    .B1(_11396_),
    .X(_11403_));
 sky130_fd_sc_hd__nand3_2 _21546_ (.A(_11402_),
    .B(_11396_),
    .C(_11400_),
    .Y(_11404_));
 sky130_fd_sc_hd__o22ai_4 _21547_ (.A1(_10897_),
    .A2(_11395_),
    .B1(_11399_),
    .B2(_11401_),
    .Y(_11405_));
 sky130_fd_sc_hd__and3_1 _21548_ (.A(_11405_),
    .B(_08714_),
    .C(_11404_),
    .X(_11406_));
 sky130_fd_sc_hd__nand3_1 _21549_ (.A(_11405_),
    .B(_08714_),
    .C(_11404_),
    .Y(_11407_));
 sky130_fd_sc_hd__a31oi_4 _21550_ (.A1(_11405_),
    .A2(_08714_),
    .A3(_11404_),
    .B1(_11393_),
    .Y(_11409_));
 sky130_fd_sc_hd__o211a_2 _21551_ (.A1(_06989_),
    .A2(net375),
    .B1(_11394_),
    .C1(_11407_),
    .X(_11410_));
 sky130_fd_sc_hd__a311o_1 _21552_ (.A1(_11405_),
    .A2(_08714_),
    .A3(_11404_),
    .B1(_11393_),
    .C1(_07044_),
    .X(_11411_));
 sky130_fd_sc_hd__a21oi_1 _21553_ (.A1(_11394_),
    .A2(_11407_),
    .B1(_07033_),
    .Y(_11412_));
 sky130_fd_sc_hd__a22o_1 _21554_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_11394_),
    .B2(_11407_),
    .X(_11413_));
 sky130_fd_sc_hd__o21ai_1 _21555_ (.A1(_10906_),
    .A2(_10913_),
    .B1(_11413_),
    .Y(_11414_));
 sky130_fd_sc_hd__o21ai_1 _21556_ (.A1(_11410_),
    .A2(_11412_),
    .B1(_10961_),
    .Y(_11415_));
 sky130_fd_sc_hd__nand3_1 _21557_ (.A(_11413_),
    .B(_10961_),
    .C(_11411_),
    .Y(_11416_));
 sky130_fd_sc_hd__o22ai_1 _21558_ (.A1(_10906_),
    .A2(_10913_),
    .B1(_11410_),
    .B2(_11412_),
    .Y(_11417_));
 sky130_fd_sc_hd__o211ai_2 _21559_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_11416_),
    .C1(_11417_),
    .Y(_11418_));
 sky130_fd_sc_hd__or4_1 _21560_ (.A(_09120_),
    .B(_09121_),
    .C(_11393_),
    .D(_11406_),
    .X(_11420_));
 sky130_fd_sc_hd__o211ai_2 _21561_ (.A1(_11414_),
    .A2(_11410_),
    .B1(_09125_),
    .C1(_11415_),
    .Y(_11421_));
 sky130_fd_sc_hd__nand2_1 _21562_ (.A(_11418_),
    .B(_11420_),
    .Y(_11422_));
 sky130_fd_sc_hd__or3_2 _21563_ (.A(_09553_),
    .B(net155),
    .C(_11422_),
    .X(_11423_));
 sky130_fd_sc_hd__o311a_2 _21564_ (.A1(_09125_),
    .A2(_11393_),
    .A3(_11406_),
    .B1(_11418_),
    .C1(_06343_),
    .X(_11424_));
 sky130_fd_sc_hd__o211ai_1 _21565_ (.A1(net394),
    .A2(_06267_),
    .B1(_11418_),
    .C1(_11420_),
    .Y(_11425_));
 sky130_fd_sc_hd__o221ai_4 _21566_ (.A1(net381),
    .A2(_06310_),
    .B1(_09125_),
    .B2(_11409_),
    .C1(_11421_),
    .Y(_11426_));
 sky130_fd_sc_hd__a31oi_2 _21567_ (.A1(_10917_),
    .A2(_10918_),
    .A3(_10921_),
    .B1(_10922_),
    .Y(_11427_));
 sky130_fd_sc_hd__a21o_1 _21568_ (.A1(_11425_),
    .A2(_11426_),
    .B1(_11427_),
    .X(_11428_));
 sky130_fd_sc_hd__a21boi_2 _21569_ (.A1(_11422_),
    .A2(_06332_),
    .B1_N(_11427_),
    .Y(_11429_));
 sky130_fd_sc_hd__nand2_1 _21570_ (.A(_11426_),
    .B(_11427_),
    .Y(_11431_));
 sky130_fd_sc_hd__o221ai_4 _21571_ (.A1(_09553_),
    .A2(net155),
    .B1(_11424_),
    .B2(_11431_),
    .C1(_11428_),
    .Y(_11432_));
 sky130_fd_sc_hd__o211ai_1 _21572_ (.A1(_05556_),
    .A2(_10929_),
    .B1(_10927_),
    .C1(_10925_),
    .Y(_11433_));
 sky130_fd_sc_hd__a21oi_1 _21573_ (.A1(_10931_),
    .A2(_11433_),
    .B1(_05851_),
    .Y(_11434_));
 sky130_fd_sc_hd__a22o_1 _21574_ (.A1(net395),
    .A2(_05796_),
    .B1(_10931_),
    .B2(_11433_),
    .X(_11435_));
 sky130_fd_sc_hd__and3_1 _21575_ (.A(_11433_),
    .B(_05851_),
    .C(_10931_),
    .X(_11436_));
 sky130_fd_sc_hd__a211o_1 _21576_ (.A1(_09572_),
    .A2(_09574_),
    .B1(_11434_),
    .C1(_11436_),
    .X(_11437_));
 sky130_fd_sc_hd__a21oi_2 _21577_ (.A1(_11423_),
    .A2(_11432_),
    .B1(_11437_),
    .Y(_11438_));
 sky130_fd_sc_hd__o311a_2 _21578_ (.A1(_09578_),
    .A2(_11434_),
    .A3(_11436_),
    .B1(_11423_),
    .C1(_11432_),
    .X(_11439_));
 sky130_fd_sc_hd__nor2_1 _21579_ (.A(_11438_),
    .B(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__o21ai_4 _21580_ (.A1(_10471_),
    .A2(_10940_),
    .B1(_10939_),
    .Y(_11442_));
 sky130_fd_sc_hd__o21ai_1 _21581_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_11442_),
    .Y(_11443_));
 sky130_fd_sc_hd__a21o_1 _21582_ (.A1(_05512_),
    .A2(net396),
    .B1(_11442_),
    .X(_11444_));
 sky130_fd_sc_hd__o221ai_4 _21583_ (.A1(_10474_),
    .A2(net138),
    .B1(_11442_),
    .B2(_05556_),
    .C1(_11443_),
    .Y(_11445_));
 sky130_fd_sc_hd__o21ai_2 _21584_ (.A1(_11438_),
    .A2(_11439_),
    .B1(_11445_),
    .Y(_11446_));
 sky130_fd_sc_hd__o31ai_4 _21585_ (.A1(_11438_),
    .A2(_11439_),
    .A3(_11445_),
    .B1(_11446_),
    .Y(_11447_));
 sky130_fd_sc_hd__o311a_1 _21586_ (.A1(_11438_),
    .A2(_11439_),
    .A3(_11445_),
    .B1(_05239_),
    .C1(_11446_),
    .X(_11448_));
 sky130_fd_sc_hd__o21a_1 _21587_ (.A1(net407),
    .A2(_05218_),
    .B1(_11447_),
    .X(_11449_));
 sky130_fd_sc_hd__a21oi_2 _21588_ (.A1(_05250_),
    .A2(_11447_),
    .B1(_10945_),
    .Y(_11450_));
 sky130_fd_sc_hd__o31a_1 _21589_ (.A1(net407),
    .A2(_05218_),
    .A3(_11447_),
    .B1(_11450_),
    .X(_11451_));
 sky130_fd_sc_hd__o2bb2a_1 _21590_ (.A1_N(net1),
    .A2_N(_10944_),
    .B1(_11448_),
    .B2(_11449_),
    .X(_11453_));
 sky130_fd_sc_hd__o22a_1 _21591_ (.A1(_10949_),
    .A2(net136),
    .B1(_11451_),
    .B2(_11453_),
    .X(_11454_));
 sky130_fd_sc_hd__a31o_1 _21592_ (.A1(_10950_),
    .A2(_10952_),
    .A3(_11447_),
    .B1(_11454_),
    .X(_11455_));
 sky130_fd_sc_hd__a311oi_4 _21593_ (.A1(_10950_),
    .A2(_10952_),
    .A3(_11447_),
    .B1(_03289_),
    .C1(_11454_),
    .Y(_11456_));
 sky130_fd_sc_hd__and2_1 _21594_ (.A(_03289_),
    .B(_11455_),
    .X(_11457_));
 sky130_fd_sc_hd__or3_1 _21595_ (.A(net53),
    .B(net54),
    .C(_10473_),
    .X(_11458_));
 sky130_fd_sc_hd__and3b_4 _21596_ (.A_N(net56),
    .B(_11458_),
    .C(net57),
    .X(_11459_));
 sky130_fd_sc_hd__clkinv_4 _21597_ (.A(_11459_),
    .Y(_11460_));
 sky130_fd_sc_hd__a21boi_4 _21598_ (.A1(_11458_),
    .A2(net57),
    .B1_N(net56),
    .Y(_11461_));
 sky130_fd_sc_hd__clkinv_4 _21599_ (.A(_11461_),
    .Y(_11462_));
 sky130_fd_sc_hd__nor2_8 _21600_ (.A(_11459_),
    .B(_11461_),
    .Y(_11464_));
 sky130_fd_sc_hd__nand2_8 _21601_ (.A(_11460_),
    .B(_11462_),
    .Y(_11465_));
 sky130_fd_sc_hd__a311o_1 _21602_ (.A1(_10950_),
    .A2(_10952_),
    .A3(_11447_),
    .B1(_11465_),
    .C1(_11454_),
    .X(_11466_));
 sky130_fd_sc_hd__o31a_1 _21603_ (.A1(_11456_),
    .A2(_11457_),
    .A3(_11464_),
    .B1(_11466_),
    .X(_11467_));
 sky130_fd_sc_hd__xnor2_1 _21604_ (.A(_10960_),
    .B(_11467_),
    .Y(net88));
 sky130_fd_sc_hd__nand3_2 _21605_ (.A(_10483_),
    .B(_10956_),
    .C(_11467_),
    .Y(_11468_));
 sky130_fd_sc_hd__or4_4 _21606_ (.A(_03399_),
    .B(net21),
    .C(net22),
    .D(_10020_),
    .X(_11469_));
 sky130_fd_sc_hd__nor2_8 _21607_ (.A(net24),
    .B(_11469_),
    .Y(_11470_));
 sky130_fd_sc_hd__or4_4 _21608_ (.A(_03399_),
    .B(net22),
    .C(net24),
    .D(_10485_),
    .X(_11471_));
 sky130_fd_sc_hd__or4_2 _21609_ (.A(_03178_),
    .B(_03399_),
    .C(net24),
    .D(_10962_),
    .X(_11472_));
 sky130_fd_sc_hd__or4_1 _21610_ (.A(_03178_),
    .B(net24),
    .C(net405),
    .D(_11469_),
    .X(_11474_));
 sky130_fd_sc_hd__a22o_1 _21611_ (.A1(_10966_),
    .A2(_10968_),
    .B1(_11470_),
    .B2(net33),
    .X(_11475_));
 sky130_fd_sc_hd__a22oi_4 _21612_ (.A1(_10970_),
    .A2(_11472_),
    .B1(_10981_),
    .B2(_10975_),
    .Y(_11476_));
 sky130_fd_sc_hd__o21ai_2 _21613_ (.A1(_11475_),
    .A2(_10979_),
    .B1(net405),
    .Y(_11477_));
 sky130_fd_sc_hd__o22ai_4 _21614_ (.A1(net405),
    .A2(_11472_),
    .B1(_11477_),
    .B2(_11476_),
    .Y(_11478_));
 sky130_fd_sc_hd__or3b_1 _21615_ (.A(_05348_),
    .B(net401),
    .C_N(_11478_),
    .X(_11479_));
 sky130_fd_sc_hd__o21ai_2 _21616_ (.A1(_10487_),
    .A2(_10488_),
    .B1(_11478_),
    .Y(_11480_));
 sky130_fd_sc_hd__o211ai_2 _21617_ (.A1(_11477_),
    .A2(_11476_),
    .B1(_11474_),
    .C1(net150),
    .Y(_11481_));
 sky130_fd_sc_hd__and2_1 _21618_ (.A(_11480_),
    .B(_11481_),
    .X(_11482_));
 sky130_fd_sc_hd__nand2_1 _21619_ (.A(_11480_),
    .B(_11481_),
    .Y(_11483_));
 sky130_fd_sc_hd__o31ai_1 _21620_ (.A1(_10989_),
    .A2(_10998_),
    .A3(_11003_),
    .B1(_10988_),
    .Y(_11485_));
 sky130_fd_sc_hd__o21bai_4 _21621_ (.A1(_10987_),
    .A2(_11006_),
    .B1_N(_11483_),
    .Y(_11486_));
 sky130_fd_sc_hd__a21oi_1 _21622_ (.A1(_11480_),
    .A2(_11481_),
    .B1(_10987_),
    .Y(_11487_));
 sky130_fd_sc_hd__a22oi_4 _21623_ (.A1(_05359_),
    .A2(_05381_),
    .B1(_11007_),
    .B2(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__nand2_1 _21624_ (.A(_11486_),
    .B(_11488_),
    .Y(_11489_));
 sky130_fd_sc_hd__a22oi_4 _21625_ (.A1(_05392_),
    .A2(_11478_),
    .B1(_11486_),
    .B2(_11488_),
    .Y(_11490_));
 sky130_fd_sc_hd__a22o_1 _21626_ (.A1(_05392_),
    .A2(_11478_),
    .B1(_11486_),
    .B2(_11488_),
    .X(_11491_));
 sky130_fd_sc_hd__or3_2 _21627_ (.A(_05676_),
    .B(_05698_),
    .C(_11490_),
    .X(_11492_));
 sky130_fd_sc_hd__a21oi_1 _21628_ (.A1(_11479_),
    .A2(_11489_),
    .B1(_10026_),
    .Y(_11493_));
 sky130_fd_sc_hd__o21ai_2 _21629_ (.A1(_10021_),
    .A2(_10022_),
    .B1(_11491_),
    .Y(_11494_));
 sky130_fd_sc_hd__and3_1 _21630_ (.A(_11489_),
    .B(_10026_),
    .C(_11479_),
    .X(_11496_));
 sky130_fd_sc_hd__o21ai_1 _21631_ (.A1(_10023_),
    .A2(_10024_),
    .B1(_11490_),
    .Y(_11497_));
 sky130_fd_sc_hd__nor2_1 _21632_ (.A(_11493_),
    .B(_11496_),
    .Y(_11498_));
 sky130_fd_sc_hd__nand2_2 _21633_ (.A(_11494_),
    .B(_11497_),
    .Y(_11499_));
 sky130_fd_sc_hd__a21oi_1 _21634_ (.A1(net175),
    .A2(_10055_),
    .B1(_09630_),
    .Y(_11500_));
 sky130_fd_sc_hd__and3_1 _21635_ (.A(_10060_),
    .B(_10062_),
    .C(_09629_),
    .X(_11501_));
 sky130_fd_sc_hd__nand4_2 _21636_ (.A(_10527_),
    .B(_11500_),
    .C(_10528_),
    .D(_10062_),
    .Y(_11502_));
 sky130_fd_sc_hd__nand4_1 _21637_ (.A(_11501_),
    .B(_11018_),
    .C(_10528_),
    .D(_10527_),
    .Y(_11503_));
 sky130_fd_sc_hd__o32ai_4 _21638_ (.A1(net172),
    .A2(_11009_),
    .A3(_11010_),
    .B1(_11502_),
    .B2(_11017_),
    .Y(_11504_));
 sky130_fd_sc_hd__a31oi_4 _21639_ (.A1(_11020_),
    .A2(_11015_),
    .A3(_10528_),
    .B1(_11504_),
    .Y(_11505_));
 sky130_fd_sc_hd__a31o_1 _21640_ (.A1(_11020_),
    .A2(_11015_),
    .A3(_10528_),
    .B1(_11504_),
    .X(_11507_));
 sky130_fd_sc_hd__nor3_2 _21641_ (.A(_09641_),
    .B(_11019_),
    .C(_11503_),
    .Y(_11508_));
 sky130_fd_sc_hd__a211o_1 _21642_ (.A1(_09595_),
    .A2(_11012_),
    .B1(_09641_),
    .C1(_11503_),
    .X(_11509_));
 sky130_fd_sc_hd__a21oi_2 _21643_ (.A1(_11507_),
    .A2(_11509_),
    .B1(_11498_),
    .Y(_11510_));
 sky130_fd_sc_hd__o21ai_1 _21644_ (.A1(_11505_),
    .A2(_11508_),
    .B1(_11499_),
    .Y(_11511_));
 sky130_fd_sc_hd__nor3_1 _21645_ (.A(_11508_),
    .B(_11499_),
    .C(_11505_),
    .Y(_11512_));
 sky130_fd_sc_hd__nand3_2 _21646_ (.A(_11507_),
    .B(_11509_),
    .C(_11498_),
    .Y(_11513_));
 sky130_fd_sc_hd__o31ai_4 _21647_ (.A1(_11508_),
    .A2(_11499_),
    .A3(_11505_),
    .B1(net358),
    .Y(_11514_));
 sky130_fd_sc_hd__nand3_2 _21648_ (.A(_11511_),
    .B(_11513_),
    .C(net358),
    .Y(_11515_));
 sky130_fd_sc_hd__o22ai_1 _21649_ (.A1(net358),
    .A2(_11490_),
    .B1(_11510_),
    .B2(_11514_),
    .Y(_11516_));
 sky130_fd_sc_hd__and3_2 _21650_ (.A(_06804_),
    .B(_06826_),
    .C(_11516_),
    .X(_11518_));
 sky130_fd_sc_hd__a211o_1 _21651_ (.A1(_11492_),
    .A2(_11515_),
    .B1(_06793_),
    .C1(_06815_),
    .X(_11519_));
 sky130_fd_sc_hd__a2bb2oi_4 _21652_ (.A1_N(_09588_),
    .A2_N(net187),
    .B1(_11492_),
    .B2(_11515_),
    .Y(_11520_));
 sky130_fd_sc_hd__o21ai_2 _21653_ (.A1(_09588_),
    .A2(net187),
    .B1(_11516_),
    .Y(_11521_));
 sky130_fd_sc_hd__o22a_1 _21654_ (.A1(_09592_),
    .A2(_09593_),
    .B1(_11510_),
    .B2(_11514_),
    .X(_11522_));
 sky130_fd_sc_hd__o221a_1 _21655_ (.A1(net358),
    .A2(_11490_),
    .B1(_11510_),
    .B2(_11514_),
    .C1(net172),
    .X(_11523_));
 sky130_fd_sc_hd__o221ai_4 _21656_ (.A1(net358),
    .A2(_11490_),
    .B1(_11510_),
    .B2(_11514_),
    .C1(net172),
    .Y(_11524_));
 sky130_fd_sc_hd__a21oi_1 _21657_ (.A1(_11492_),
    .A2(_11522_),
    .B1(_11520_),
    .Y(_11525_));
 sky130_fd_sc_hd__nand2_1 _21658_ (.A(_11521_),
    .B(_11524_),
    .Y(_11526_));
 sky130_fd_sc_hd__o211ai_2 _21659_ (.A1(_10547_),
    .A2(_10548_),
    .B1(_11029_),
    .C1(_10543_),
    .Y(_11527_));
 sky130_fd_sc_hd__o2111ai_4 _21660_ (.A1(net173),
    .A2(_11025_),
    .B1(_11521_),
    .C1(_11524_),
    .D1(_11527_),
    .Y(_11529_));
 sky130_fd_sc_hd__o211ai_4 _21661_ (.A1(_11520_),
    .A2(_11523_),
    .B1(_11029_),
    .C1(_11033_),
    .Y(_11530_));
 sky130_fd_sc_hd__nand3_1 _21662_ (.A(_11530_),
    .B(net357),
    .C(_11529_),
    .Y(_11531_));
 sky130_fd_sc_hd__a31oi_4 _21663_ (.A1(_11530_),
    .A2(net357),
    .A3(_11529_),
    .B1(_11518_),
    .Y(_11532_));
 sky130_fd_sc_hd__a2bb2oi_2 _21664_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_11519_),
    .B2(_11531_),
    .Y(_11533_));
 sky130_fd_sc_hd__a311oi_4 _21665_ (.A1(_11530_),
    .A2(net357),
    .A3(_11529_),
    .B1(net173),
    .C1(_11518_),
    .Y(_11534_));
 sky130_fd_sc_hd__a311o_2 _21666_ (.A1(_11530_),
    .A2(net357),
    .A3(_11529_),
    .B1(net173),
    .C1(_11518_),
    .X(_11535_));
 sky130_fd_sc_hd__nor2_1 _21667_ (.A(_11533_),
    .B(_11534_),
    .Y(_11536_));
 sky130_fd_sc_hd__o32ai_1 _21668_ (.A1(net177),
    .A2(_11026_),
    .A3(_11036_),
    .B1(_11047_),
    .B2(_11048_),
    .Y(_11537_));
 sky130_fd_sc_hd__o221ai_4 _21669_ (.A1(_11533_),
    .A2(_11534_),
    .B1(_11047_),
    .B2(_11048_),
    .C1(_11043_),
    .Y(_11538_));
 sky130_fd_sc_hd__nand2_1 _21670_ (.A(_11537_),
    .B(_11536_),
    .Y(_11540_));
 sky130_fd_sc_hd__or3_1 _21671_ (.A(net374),
    .B(_07702_),
    .C(_11532_),
    .X(_11541_));
 sky130_fd_sc_hd__nand3_4 _21672_ (.A(_11540_),
    .B(net355),
    .C(_11538_),
    .Y(_11542_));
 sky130_fd_sc_hd__o31a_1 _21673_ (.A1(net374),
    .A2(_07702_),
    .A3(_11532_),
    .B1(_11542_),
    .X(_11543_));
 sky130_fd_sc_hd__a21oi_1 _21674_ (.A1(_11541_),
    .A2(_11542_),
    .B1(net338),
    .Y(_11544_));
 sky130_fd_sc_hd__or3_2 _21675_ (.A(_08678_),
    .B(_08700_),
    .C(_11543_),
    .X(_11545_));
 sky130_fd_sc_hd__a2bb2oi_2 _21676_ (.A1_N(_08724_),
    .A2_N(_08726_),
    .B1(_11541_),
    .B2(_11542_),
    .Y(_11546_));
 sky130_fd_sc_hd__a22o_2 _21677_ (.A1(_08725_),
    .A2(_08727_),
    .B1(_11541_),
    .B2(_11542_),
    .X(_11547_));
 sky130_fd_sc_hd__o211a_2 _21678_ (.A1(net354),
    .A2(_11532_),
    .B1(net177),
    .C1(_11542_),
    .X(_11548_));
 sky130_fd_sc_hd__o211ai_4 _21679_ (.A1(net354),
    .A2(_11532_),
    .B1(net177),
    .C1(_11542_),
    .Y(_11549_));
 sky130_fd_sc_hd__a2bb2oi_1 _21680_ (.A1_N(net199),
    .A2_N(_11052_),
    .B1(_11066_),
    .B2(_11070_),
    .Y(_11551_));
 sky130_fd_sc_hd__o31ai_2 _21681_ (.A1(_11064_),
    .A2(_10591_),
    .A3(_10589_),
    .B1(_11058_),
    .Y(_11552_));
 sky130_fd_sc_hd__o22ai_4 _21682_ (.A1(net199),
    .A2(_11052_),
    .B1(_11552_),
    .B2(_11069_),
    .Y(_11553_));
 sky130_fd_sc_hd__a31oi_2 _21683_ (.A1(_11058_),
    .A2(_11066_),
    .A3(_11070_),
    .B1(_11054_),
    .Y(_11554_));
 sky130_fd_sc_hd__nand3_4 _21684_ (.A(_11553_),
    .B(_11549_),
    .C(_11547_),
    .Y(_11555_));
 sky130_fd_sc_hd__o211ai_4 _21685_ (.A1(_11546_),
    .A2(_11548_),
    .B1(_11055_),
    .C1(_11076_),
    .Y(_11556_));
 sky130_fd_sc_hd__nand3_2 _21686_ (.A(_11555_),
    .B(_11556_),
    .C(net338),
    .Y(_11557_));
 sky130_fd_sc_hd__o311a_1 _21687_ (.A1(net374),
    .A2(_07702_),
    .A3(_11532_),
    .B1(_11542_),
    .C1(_08732_),
    .X(_11558_));
 sky130_fd_sc_hd__a22oi_2 _21688_ (.A1(_08689_),
    .A2(_08711_),
    .B1(_11555_),
    .B2(_11556_),
    .Y(_11559_));
 sky130_fd_sc_hd__o31a_1 _21689_ (.A1(_08678_),
    .A2(_08700_),
    .A3(_11543_),
    .B1(_11557_),
    .X(_11560_));
 sky130_fd_sc_hd__a31o_2 _21690_ (.A1(_11555_),
    .A2(_11556_),
    .A3(net338),
    .B1(_11544_),
    .X(_11562_));
 sky130_fd_sc_hd__a2bb2oi_2 _21691_ (.A1_N(_08307_),
    .A2_N(_08309_),
    .B1(_11545_),
    .B2(_11557_),
    .Y(_11563_));
 sky130_fd_sc_hd__a22o_2 _21692_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_11545_),
    .B2(_11557_),
    .X(_11564_));
 sky130_fd_sc_hd__a31oi_2 _21693_ (.A1(_11555_),
    .A2(_11556_),
    .A3(net338),
    .B1(net198),
    .Y(_11565_));
 sky130_fd_sc_hd__o221a_1 _21694_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_11543_),
    .B2(net338),
    .C1(_11557_),
    .X(_11566_));
 sky130_fd_sc_hd__a311o_2 _21695_ (.A1(_11555_),
    .A2(_11556_),
    .A3(net338),
    .B1(net198),
    .C1(_11544_),
    .X(_11567_));
 sky130_fd_sc_hd__a21oi_4 _21696_ (.A1(_11545_),
    .A2(_11565_),
    .B1(_11563_),
    .Y(_11568_));
 sky130_fd_sc_hd__o41ai_1 _21697_ (.A1(_08311_),
    .A2(_08312_),
    .A3(_11558_),
    .A4(_11559_),
    .B1(_11567_),
    .Y(_11569_));
 sky130_fd_sc_hd__nor3_1 _21698_ (.A(_10139_),
    .B(_09710_),
    .C(_10137_),
    .Y(_11570_));
 sky130_fd_sc_hd__nor3b_2 _21699_ (.A(_10599_),
    .B(_10601_),
    .C_N(_11570_),
    .Y(_11571_));
 sky130_fd_sc_hd__nand3_1 _21700_ (.A(_10600_),
    .B(_10602_),
    .C(_11570_),
    .Y(_11573_));
 sky130_fd_sc_hd__nand3_2 _21701_ (.A(_11571_),
    .B(_11091_),
    .C(_11088_),
    .Y(_11574_));
 sky130_fd_sc_hd__nand4_4 _21702_ (.A(_11571_),
    .B(_11091_),
    .C(_11088_),
    .D(_09718_),
    .Y(_11575_));
 sky130_fd_sc_hd__a21oi_1 _21703_ (.A1(_11571_),
    .A2(_11091_),
    .B1(_11087_),
    .Y(_11576_));
 sky130_fd_sc_hd__o211ai_4 _21704_ (.A1(_11573_),
    .A2(_11089_),
    .B1(_11088_),
    .C1(_11092_),
    .Y(_11577_));
 sky130_fd_sc_hd__a2bb2oi_4 _21705_ (.A1_N(_09720_),
    .A2_N(_11574_),
    .B1(_11094_),
    .B2(_11576_),
    .Y(_11578_));
 sky130_fd_sc_hd__o21ai_2 _21706_ (.A1(_09720_),
    .A2(_11574_),
    .B1(_11577_),
    .Y(_11579_));
 sky130_fd_sc_hd__a21oi_2 _21707_ (.A1(_11575_),
    .A2(_11577_),
    .B1(_11569_),
    .Y(_11580_));
 sky130_fd_sc_hd__o22ai_2 _21708_ (.A1(net351),
    .A2(_09807_),
    .B1(_11568_),
    .B2(_11579_),
    .Y(_11581_));
 sky130_fd_sc_hd__nand4_4 _21709_ (.A(_11564_),
    .B(_11567_),
    .C(_11575_),
    .D(_11577_),
    .Y(_11582_));
 sky130_fd_sc_hd__o21ai_2 _21710_ (.A1(_11563_),
    .A2(_11566_),
    .B1(_11579_),
    .Y(_11584_));
 sky130_fd_sc_hd__o221ai_4 _21711_ (.A1(net351),
    .A2(_09807_),
    .B1(_11568_),
    .B2(_11578_),
    .C1(_11582_),
    .Y(_11585_));
 sky130_fd_sc_hd__a2bb2o_2 _21712_ (.A1_N(_09763_),
    .A2_N(_09774_),
    .B1(_11545_),
    .B2(_11557_),
    .X(_11586_));
 sky130_fd_sc_hd__inv_2 _21713_ (.A(_11586_),
    .Y(_11587_));
 sky130_fd_sc_hd__a31o_1 _21714_ (.A1(_11584_),
    .A2(net335),
    .A3(_11582_),
    .B1(_11587_),
    .X(_11588_));
 sky130_fd_sc_hd__o221a_2 _21715_ (.A1(net335),
    .A2(_11562_),
    .B1(_11580_),
    .B2(_11581_),
    .C1(_11079_),
    .X(_11589_));
 sky130_fd_sc_hd__a211o_1 _21716_ (.A1(_11585_),
    .A2(_11586_),
    .B1(_11046_),
    .C1(_11057_),
    .X(_11590_));
 sky130_fd_sc_hd__o211a_1 _21717_ (.A1(_10614_),
    .A2(net224),
    .B1(_11109_),
    .C1(_11103_),
    .X(_11591_));
 sky130_fd_sc_hd__o211a_1 _21718_ (.A1(_10613_),
    .A2(net222),
    .B1(_11108_),
    .C1(_11106_),
    .X(_11592_));
 sky130_fd_sc_hd__a31oi_2 _21719_ (.A1(_10616_),
    .A2(_11106_),
    .A3(_11108_),
    .B1(_11102_),
    .Y(_11593_));
 sky130_fd_sc_hd__a311oi_4 _21720_ (.A1(_11584_),
    .A2(net335),
    .A3(_11582_),
    .B1(_11587_),
    .C1(_07936_),
    .Y(_11595_));
 sky130_fd_sc_hd__nand3_4 _21721_ (.A(_11585_),
    .B(_11586_),
    .C(_07935_),
    .Y(_11596_));
 sky130_fd_sc_hd__a21oi_1 _21722_ (.A1(_11585_),
    .A2(_11586_),
    .B1(_07935_),
    .Y(_11597_));
 sky130_fd_sc_hd__o221ai_4 _21723_ (.A1(net335),
    .A2(_11562_),
    .B1(_11580_),
    .B2(_11581_),
    .C1(_07936_),
    .Y(_11598_));
 sky130_fd_sc_hd__o211a_1 _21724_ (.A1(_11102_),
    .A2(_11592_),
    .B1(_11596_),
    .C1(_11598_),
    .X(_11599_));
 sky130_fd_sc_hd__o211ai_4 _21725_ (.A1(_11102_),
    .A2(_11592_),
    .B1(_11596_),
    .C1(_11598_),
    .Y(_11600_));
 sky130_fd_sc_hd__a21boi_1 _21726_ (.A1(_11596_),
    .A2(_11598_),
    .B1_N(_11593_),
    .Y(_11601_));
 sky130_fd_sc_hd__o22ai_4 _21727_ (.A1(_11105_),
    .A2(_11591_),
    .B1(_11595_),
    .B2(_11597_),
    .Y(_11602_));
 sky130_fd_sc_hd__nand3_2 _21728_ (.A(_11602_),
    .B(net332),
    .C(_11600_),
    .Y(_11603_));
 sky130_fd_sc_hd__o22ai_2 _21729_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_11599_),
    .B2(_11601_),
    .Y(_11604_));
 sky130_fd_sc_hd__a31oi_4 _21730_ (.A1(_11602_),
    .A2(net332),
    .A3(_11600_),
    .B1(_11589_),
    .Y(_11606_));
 sky130_fd_sc_hd__a31o_1 _21731_ (.A1(_11602_),
    .A2(net332),
    .A3(_11600_),
    .B1(_11589_),
    .X(_11607_));
 sky130_fd_sc_hd__a311oi_4 _21732_ (.A1(_11602_),
    .A2(net332),
    .A3(_11600_),
    .B1(net202),
    .C1(_11589_),
    .Y(_11608_));
 sky130_fd_sc_hd__o211ai_4 _21733_ (.A1(_07560_),
    .A2(_07562_),
    .B1(_11590_),
    .C1(_11603_),
    .Y(_11609_));
 sky130_fd_sc_hd__a2bb2oi_2 _21734_ (.A1_N(_07555_),
    .A2_N(net218),
    .B1(_11590_),
    .B2(_11603_),
    .Y(_11610_));
 sky130_fd_sc_hd__o221ai_4 _21735_ (.A1(_07555_),
    .A2(net218),
    .B1(_11588_),
    .B2(net332),
    .C1(_11604_),
    .Y(_11611_));
 sky130_fd_sc_hd__nor2_1 _21736_ (.A(_11608_),
    .B(_11610_),
    .Y(_11612_));
 sky130_fd_sc_hd__o211ai_4 _21737_ (.A1(net227),
    .A2(_10626_),
    .B1(_11120_),
    .C1(_11125_),
    .Y(_11613_));
 sky130_fd_sc_hd__a31oi_1 _21738_ (.A1(_10631_),
    .A2(_11120_),
    .A3(_11125_),
    .B1(_11121_),
    .Y(_11614_));
 sky130_fd_sc_hd__o21ai_1 _21739_ (.A1(net222),
    .A2(_11118_),
    .B1(_11613_),
    .Y(_11615_));
 sky130_fd_sc_hd__o2111ai_1 _21740_ (.A1(_11124_),
    .A2(_11126_),
    .B1(_11609_),
    .C1(_11611_),
    .D1(_11120_),
    .Y(_11617_));
 sky130_fd_sc_hd__o21ai_1 _21741_ (.A1(_11608_),
    .A2(_11610_),
    .B1(_11614_),
    .Y(_11618_));
 sky130_fd_sc_hd__o211ai_1 _21742_ (.A1(net329),
    .A2(net327),
    .B1(_11617_),
    .C1(_11618_),
    .Y(_11619_));
 sky130_fd_sc_hd__or3_1 _21743_ (.A(net329),
    .B(net327),
    .C(_11606_),
    .X(_11620_));
 sky130_fd_sc_hd__o21ai_1 _21744_ (.A1(_11608_),
    .A2(_11610_),
    .B1(_11615_),
    .Y(_11621_));
 sky130_fd_sc_hd__o221ai_4 _21745_ (.A1(_11118_),
    .A2(net222),
    .B1(_07564_),
    .B2(_11606_),
    .C1(_11613_),
    .Y(_11622_));
 sky130_fd_sc_hd__o221ai_4 _21746_ (.A1(net329),
    .A2(net327),
    .B1(_11608_),
    .B2(_11622_),
    .C1(_11621_),
    .Y(_11623_));
 sky130_fd_sc_hd__o31a_4 _21747_ (.A1(net329),
    .A2(net327),
    .A3(_11606_),
    .B1(_11623_),
    .X(_11624_));
 sky130_fd_sc_hd__inv_2 _21748_ (.A(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__or3_2 _21749_ (.A(_00011_),
    .B(net323),
    .C(_11624_),
    .X(_11626_));
 sky130_fd_sc_hd__o211ai_2 _21750_ (.A1(_11607_),
    .A2(net311),
    .B1(net222),
    .C1(_11619_),
    .Y(_11628_));
 sky130_fd_sc_hd__nand3_2 _21751_ (.A(_11623_),
    .B(net224),
    .C(_11620_),
    .Y(_11629_));
 sky130_fd_sc_hd__nand2_4 _21752_ (.A(_11628_),
    .B(_11629_),
    .Y(_11630_));
 sky130_fd_sc_hd__o211ai_4 _21753_ (.A1(_11138_),
    .A2(_11132_),
    .B1(_11148_),
    .C1(_11146_),
    .Y(_11631_));
 sky130_fd_sc_hd__a31oi_4 _21754_ (.A1(_11139_),
    .A2(_11146_),
    .A3(_11148_),
    .B1(_11135_),
    .Y(_11632_));
 sky130_fd_sc_hd__nand3_1 _21755_ (.A(_11136_),
    .B(_11630_),
    .C(_11631_),
    .Y(_11633_));
 sky130_fd_sc_hd__a21o_2 _21756_ (.A1(_11136_),
    .A2(_11631_),
    .B1(_11630_),
    .X(_11634_));
 sky130_fd_sc_hd__a31oi_4 _21757_ (.A1(_11136_),
    .A2(_11630_),
    .A3(_11631_),
    .B1(_00066_),
    .Y(_11635_));
 sky130_fd_sc_hd__o211ai_4 _21758_ (.A1(_11630_),
    .A2(_11632_),
    .B1(net308),
    .C1(_11633_),
    .Y(_11636_));
 sky130_fd_sc_hd__a22oi_4 _21759_ (.A1(_00066_),
    .A2(_11625_),
    .B1(_11635_),
    .B2(_11634_),
    .Y(_11637_));
 sky130_fd_sc_hd__o21ai_4 _21760_ (.A1(net307),
    .A2(_11624_),
    .B1(_11636_),
    .Y(_11639_));
 sky130_fd_sc_hd__a2bb2oi_1 _21761_ (.A1_N(_06914_),
    .A2_N(_06916_),
    .B1(_11626_),
    .B2(_11636_),
    .Y(_11640_));
 sky130_fd_sc_hd__a22o_1 _21762_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_11626_),
    .B2(_11636_),
    .X(_11641_));
 sky130_fd_sc_hd__a21oi_1 _21763_ (.A1(_11635_),
    .A2(_11634_),
    .B1(net225),
    .Y(_11642_));
 sky130_fd_sc_hd__o211a_1 _21764_ (.A1(net307),
    .A2(_11624_),
    .B1(net227),
    .C1(_11636_),
    .X(_11643_));
 sky130_fd_sc_hd__o211ai_2 _21765_ (.A1(net307),
    .A2(_11624_),
    .B1(net227),
    .C1(_11636_),
    .Y(_11644_));
 sky130_fd_sc_hd__a21oi_2 _21766_ (.A1(_11642_),
    .A2(_11626_),
    .B1(_11640_),
    .Y(_11645_));
 sky130_fd_sc_hd__nand2_1 _21767_ (.A(_11641_),
    .B(_11644_),
    .Y(_11646_));
 sky130_fd_sc_hd__and4_1 _21768_ (.A(_09778_),
    .B(_09779_),
    .C(_10207_),
    .D(_10209_),
    .X(_11647_));
 sky130_fd_sc_hd__nand4_1 _21769_ (.A(_09778_),
    .B(_09779_),
    .C(_10207_),
    .D(_10209_),
    .Y(_11648_));
 sky130_fd_sc_hd__a211oi_2 _21770_ (.A1(_10654_),
    .A2(_10672_),
    .B1(_11648_),
    .C1(_10676_),
    .Y(_11650_));
 sky130_fd_sc_hd__nand3_2 _21771_ (.A(_11162_),
    .B(_11647_),
    .C(_10678_),
    .Y(_11651_));
 sky130_fd_sc_hd__a21oi_1 _21772_ (.A1(_11650_),
    .A2(_11162_),
    .B1(_11163_),
    .Y(_11652_));
 sky130_fd_sc_hd__o211a_1 _21773_ (.A1(_11168_),
    .A2(_11161_),
    .B1(_11164_),
    .C1(_11651_),
    .X(_11653_));
 sky130_fd_sc_hd__o211ai_4 _21774_ (.A1(_11168_),
    .A2(_11161_),
    .B1(_11164_),
    .C1(_11651_),
    .Y(_11654_));
 sky130_fd_sc_hd__o2111a_1 _21775_ (.A1(_09784_),
    .A2(_09788_),
    .B1(_10675_),
    .C1(_11647_),
    .D1(_10677_),
    .X(_11655_));
 sky130_fd_sc_hd__nand3_1 _21776_ (.A(_11650_),
    .B(_11164_),
    .C(_09789_),
    .Y(_11656_));
 sky130_fd_sc_hd__nand4_4 _21777_ (.A(_11650_),
    .B(_11164_),
    .C(_11162_),
    .D(_09789_),
    .Y(_11657_));
 sky130_fd_sc_hd__a2bb2oi_1 _21778_ (.A1_N(_11161_),
    .A2_N(_11656_),
    .B1(_11170_),
    .B2(_11652_),
    .Y(_11658_));
 sky130_fd_sc_hd__a31o_1 _21779_ (.A1(_11162_),
    .A2(_11164_),
    .A3(_11655_),
    .B1(_11653_),
    .X(_11659_));
 sky130_fd_sc_hd__a21oi_2 _21780_ (.A1(_11654_),
    .A2(_11657_),
    .B1(_11646_),
    .Y(_11661_));
 sky130_fd_sc_hd__o211ai_1 _21781_ (.A1(_11640_),
    .A2(_11643_),
    .B1(_11654_),
    .C1(_11657_),
    .Y(_11662_));
 sky130_fd_sc_hd__o21ai_2 _21782_ (.A1(net304),
    .A2(_01951_),
    .B1(_11662_),
    .Y(_11663_));
 sky130_fd_sc_hd__nand3_2 _21783_ (.A(_11645_),
    .B(_11654_),
    .C(_11657_),
    .Y(_11664_));
 sky130_fd_sc_hd__a22o_1 _21784_ (.A1(_11641_),
    .A2(_11644_),
    .B1(_11654_),
    .B2(_11657_),
    .X(_11665_));
 sky130_fd_sc_hd__o221ai_4 _21785_ (.A1(net304),
    .A2(_01951_),
    .B1(_11645_),
    .B2(_11658_),
    .C1(_11664_),
    .Y(_11666_));
 sky130_fd_sc_hd__a211o_2 _21786_ (.A1(_11626_),
    .A2(_11636_),
    .B1(net304),
    .C1(_01951_),
    .X(_11667_));
 sky130_fd_sc_hd__inv_2 _21787_ (.A(_11667_),
    .Y(_11668_));
 sky130_fd_sc_hd__o221a_2 _21788_ (.A1(net279),
    .A2(_11639_),
    .B1(_11661_),
    .B2(_11663_),
    .C1(_04040_),
    .X(_11669_));
 sky130_fd_sc_hd__a211o_2 _21789_ (.A1(_11666_),
    .A2(_11667_),
    .B1(net302),
    .C1(_04019_),
    .X(_11670_));
 sky130_fd_sc_hd__a311oi_4 _21790_ (.A1(_11665_),
    .A2(net279),
    .A3(_11664_),
    .B1(_11668_),
    .C1(net232),
    .Y(_11672_));
 sky130_fd_sc_hd__nand3_4 _21791_ (.A(_11666_),
    .B(_11667_),
    .C(net234),
    .Y(_11673_));
 sky130_fd_sc_hd__a22oi_1 _21792_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_11666_),
    .B2(_11667_),
    .Y(_11674_));
 sky130_fd_sc_hd__o221ai_4 _21793_ (.A1(net279),
    .A2(_11639_),
    .B1(_11661_),
    .B2(_11663_),
    .C1(net232),
    .Y(_11675_));
 sky130_fd_sc_hd__a21oi_2 _21794_ (.A1(_10693_),
    .A2(_11173_),
    .B1(_11180_),
    .Y(_11676_));
 sky130_fd_sc_hd__a31o_1 _21795_ (.A1(_10693_),
    .A2(_11173_),
    .A3(_11179_),
    .B1(_11180_),
    .X(_11677_));
 sky130_fd_sc_hd__a31oi_2 _21796_ (.A1(_10693_),
    .A2(_11173_),
    .A3(_11179_),
    .B1(_11180_),
    .Y(_11678_));
 sky130_fd_sc_hd__o2bb2ai_4 _21797_ (.A1_N(_11673_),
    .A2_N(_11675_),
    .B1(_11676_),
    .B2(_11178_),
    .Y(_11679_));
 sky130_fd_sc_hd__nand3_4 _21798_ (.A(_11677_),
    .B(_11675_),
    .C(_11673_),
    .Y(_11680_));
 sky130_fd_sc_hd__nand3_2 _21799_ (.A(_11679_),
    .B(_11680_),
    .C(net277),
    .Y(_11681_));
 sky130_fd_sc_hd__a31oi_4 _21800_ (.A1(_11679_),
    .A2(_11680_),
    .A3(net277),
    .B1(_11669_),
    .Y(_11683_));
 sky130_fd_sc_hd__inv_2 _21801_ (.A(_11683_),
    .Y(_11684_));
 sky130_fd_sc_hd__o221ai_4 _21802_ (.A1(net262),
    .A2(_10705_),
    .B1(net254),
    .B2(_11191_),
    .C1(_11198_),
    .Y(_11685_));
 sky130_fd_sc_hd__o221ai_2 _21803_ (.A1(net261),
    .A2(_10704_),
    .B1(_11190_),
    .B2(net253),
    .C1(_11197_),
    .Y(_11686_));
 sky130_fd_sc_hd__a311oi_4 _21804_ (.A1(_11679_),
    .A2(_11680_),
    .A3(net277),
    .B1(net251),
    .C1(_11669_),
    .Y(_11687_));
 sky130_fd_sc_hd__nand3_2 _21805_ (.A(_11681_),
    .B(_06314_),
    .C(_11670_),
    .Y(_11688_));
 sky130_fd_sc_hd__a2bb2oi_4 _21806_ (.A1_N(_06305_),
    .A2_N(_06307_),
    .B1(_11670_),
    .B2(_11681_),
    .Y(_11689_));
 sky130_fd_sc_hd__a22o_1 _21807_ (.A1(_06306_),
    .A2(_06308_),
    .B1(_11670_),
    .B2(_11681_),
    .X(_11690_));
 sky130_fd_sc_hd__o2111ai_1 _21808_ (.A1(net254),
    .A2(_11191_),
    .B1(_11686_),
    .C1(_11688_),
    .D1(_11690_),
    .Y(_11691_));
 sky130_fd_sc_hd__o2bb2ai_1 _21809_ (.A1_N(_11195_),
    .A2_N(_11686_),
    .B1(_11687_),
    .B2(_11689_),
    .Y(_11692_));
 sky130_fd_sc_hd__nand3_2 _21810_ (.A(_11691_),
    .B(_11692_),
    .C(net272),
    .Y(_11694_));
 sky130_fd_sc_hd__or3_1 _21811_ (.A(net296),
    .B(_05232_),
    .C(_11683_),
    .X(_11695_));
 sky130_fd_sc_hd__o221ai_4 _21812_ (.A1(_11190_),
    .A2(net253),
    .B1(_06314_),
    .B2(_11683_),
    .C1(_11685_),
    .Y(_11696_));
 sky130_fd_sc_hd__o2bb2ai_1 _21813_ (.A1_N(_11194_),
    .A2_N(_11685_),
    .B1(_11687_),
    .B2(_11689_),
    .Y(_11697_));
 sky130_fd_sc_hd__o221ai_4 _21814_ (.A1(_05231_),
    .A2(_05232_),
    .B1(_11687_),
    .B2(_11696_),
    .C1(_11697_),
    .Y(_11698_));
 sky130_fd_sc_hd__o31a_2 _21815_ (.A1(net296),
    .A2(_05232_),
    .A3(_11683_),
    .B1(_11698_),
    .X(_11699_));
 sky130_fd_sc_hd__o211a_1 _21816_ (.A1(_11684_),
    .A2(net272),
    .B1(net253),
    .C1(_11694_),
    .X(_11700_));
 sky130_fd_sc_hd__o211ai_4 _21817_ (.A1(_11684_),
    .A2(net272),
    .B1(net253),
    .C1(_11694_),
    .Y(_11701_));
 sky130_fd_sc_hd__o221a_1 _21818_ (.A1(_06011_),
    .A2(_06012_),
    .B1(_11683_),
    .B2(net272),
    .C1(_11698_),
    .X(_11702_));
 sky130_fd_sc_hd__nand3_2 _21819_ (.A(_11698_),
    .B(net254),
    .C(_11695_),
    .Y(_11703_));
 sky130_fd_sc_hd__nand2_1 _21820_ (.A(_11701_),
    .B(_11703_),
    .Y(_11705_));
 sky130_fd_sc_hd__o2bb2ai_1 _21821_ (.A1_N(_11222_),
    .A2_N(_11223_),
    .B1(net262),
    .B2(_11209_),
    .Y(_11706_));
 sky130_fd_sc_hd__a31oi_2 _21822_ (.A1(_11213_),
    .A2(_11222_),
    .A3(_11223_),
    .B1(_11211_),
    .Y(_11707_));
 sky130_fd_sc_hd__a221oi_4 _21823_ (.A1(_11701_),
    .A2(_11703_),
    .B1(_11227_),
    .B2(_11222_),
    .C1(_11211_),
    .Y(_11708_));
 sky130_fd_sc_hd__o211ai_1 _21824_ (.A1(net262),
    .A2(_11209_),
    .B1(_11228_),
    .C1(_11705_),
    .Y(_11709_));
 sky130_fd_sc_hd__o2111ai_1 _21825_ (.A1(net261),
    .A2(_11208_),
    .B1(_11701_),
    .C1(_11703_),
    .D1(_11706_),
    .Y(_11710_));
 sky130_fd_sc_hd__o22ai_4 _21826_ (.A1(net270),
    .A2(_05483_),
    .B1(_11705_),
    .B2(_11707_),
    .Y(_11711_));
 sky130_fd_sc_hd__o211ai_2 _21827_ (.A1(_05481_),
    .A2(_05483_),
    .B1(_11709_),
    .C1(_11710_),
    .Y(_11712_));
 sky130_fd_sc_hd__or3_2 _21828_ (.A(net270),
    .B(_05483_),
    .C(_11699_),
    .X(_11713_));
 sky130_fd_sc_hd__inv_2 _21829_ (.A(_11713_),
    .Y(_11714_));
 sky130_fd_sc_hd__o22ai_4 _21830_ (.A1(net245),
    .A2(_11699_),
    .B1(_11708_),
    .B2(_11711_),
    .Y(_11716_));
 sky130_fd_sc_hd__o221a_1 _21831_ (.A1(net245),
    .A2(_11699_),
    .B1(_11708_),
    .B2(_11711_),
    .C1(_05754_),
    .X(_11717_));
 sky130_fd_sc_hd__a22oi_4 _21832_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_11712_),
    .B2(_11713_),
    .Y(_11718_));
 sky130_fd_sc_hd__o21ai_4 _21833_ (.A1(_05760_),
    .A2(_05762_),
    .B1(_11716_),
    .Y(_11719_));
 sky130_fd_sc_hd__o21ai_4 _21834_ (.A1(_11708_),
    .A2(_11711_),
    .B1(net263),
    .Y(_11720_));
 sky130_fd_sc_hd__o221a_2 _21835_ (.A1(net245),
    .A2(_11699_),
    .B1(_11708_),
    .B2(_11711_),
    .C1(net262),
    .X(_11721_));
 sky130_fd_sc_hd__o221ai_4 _21836_ (.A1(net246),
    .A2(_11699_),
    .B1(_11708_),
    .B2(_11711_),
    .C1(net263),
    .Y(_11722_));
 sky130_fd_sc_hd__o21ai_2 _21837_ (.A1(net267),
    .A2(_11234_),
    .B1(_11244_),
    .Y(_11723_));
 sky130_fd_sc_hd__o22a_1 _21838_ (.A1(_11237_),
    .A2(_11231_),
    .B1(_11242_),
    .B2(_11240_),
    .X(_11724_));
 sky130_fd_sc_hd__o22ai_4 _21839_ (.A1(_11237_),
    .A2(_11231_),
    .B1(_11242_),
    .B2(_11240_),
    .Y(_11725_));
 sky130_fd_sc_hd__o211ai_4 _21840_ (.A1(_11720_),
    .A2(_11714_),
    .B1(_11719_),
    .C1(_11725_),
    .Y(_11727_));
 sky130_fd_sc_hd__o21ai_2 _21841_ (.A1(_11718_),
    .A2(_11721_),
    .B1(_11724_),
    .Y(_11728_));
 sky130_fd_sc_hd__o211ai_2 _21842_ (.A1(net266),
    .A2(_05751_),
    .B1(_11727_),
    .C1(_11728_),
    .Y(_11729_));
 sky130_fd_sc_hd__a211o_1 _21843_ (.A1(_11712_),
    .A2(_11713_),
    .B1(net266),
    .C1(_05751_),
    .X(_11730_));
 sky130_fd_sc_hd__o21ai_1 _21844_ (.A1(_11718_),
    .A2(_11721_),
    .B1(_11725_),
    .Y(_11731_));
 sky130_fd_sc_hd__nand4_1 _21845_ (.A(_11239_),
    .B(_11719_),
    .C(_11722_),
    .D(_11723_),
    .Y(_11732_));
 sky130_fd_sc_hd__nand3_1 _21846_ (.A(_11731_),
    .B(_11732_),
    .C(net242),
    .Y(_11733_));
 sky130_fd_sc_hd__a31oi_4 _21847_ (.A1(_11728_),
    .A2(net242),
    .A3(_11727_),
    .B1(_11717_),
    .Y(_11734_));
 sky130_fd_sc_hd__inv_2 _21848_ (.A(_11734_),
    .Y(_11735_));
 sky130_fd_sc_hd__and3_1 _21849_ (.A(_11734_),
    .B(_05993_),
    .C(_05991_),
    .X(_11736_));
 sky130_fd_sc_hd__inv_2 _21850_ (.A(_11736_),
    .Y(_11738_));
 sky130_fd_sc_hd__o211a_1 _21851_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_11730_),
    .C1(_11733_),
    .X(_11739_));
 sky130_fd_sc_hd__o211ai_4 _21852_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_11730_),
    .C1(_11733_),
    .Y(_11740_));
 sky130_fd_sc_hd__o211ai_4 _21853_ (.A1(_11716_),
    .A2(net242),
    .B1(net292),
    .C1(_11729_),
    .Y(_11741_));
 sky130_fd_sc_hd__nand2_1 _21854_ (.A(_11740_),
    .B(_11741_),
    .Y(_11742_));
 sky130_fd_sc_hd__a21oi_1 _21855_ (.A1(net294),
    .A2(_11252_),
    .B1(_11257_),
    .Y(_11743_));
 sky130_fd_sc_hd__o21ai_2 _21856_ (.A1(_10766_),
    .A2(_11255_),
    .B1(_11262_),
    .Y(_11744_));
 sky130_fd_sc_hd__o21ai_1 _21857_ (.A1(_10764_),
    .A2(_11256_),
    .B1(_11260_),
    .Y(_11745_));
 sky130_fd_sc_hd__a21oi_2 _21858_ (.A1(_11260_),
    .A2(_11257_),
    .B1(_11261_),
    .Y(_11746_));
 sky130_fd_sc_hd__a22oi_1 _21859_ (.A1(_11740_),
    .A2(_11741_),
    .B1(_11744_),
    .B2(_11260_),
    .Y(_11747_));
 sky130_fd_sc_hd__o2bb2ai_1 _21860_ (.A1_N(_11740_),
    .A2_N(_11741_),
    .B1(_11743_),
    .B2(_11259_),
    .Y(_11749_));
 sky130_fd_sc_hd__a22oi_2 _21861_ (.A1(_11734_),
    .A2(net292),
    .B1(_11262_),
    .B2(_11745_),
    .Y(_11750_));
 sky130_fd_sc_hd__o2111a_1 _21862_ (.A1(net294),
    .A2(_11252_),
    .B1(_11740_),
    .C1(_11741_),
    .D1(_11744_),
    .X(_11751_));
 sky130_fd_sc_hd__o2111ai_4 _21863_ (.A1(net294),
    .A2(_11252_),
    .B1(_11740_),
    .C1(_11741_),
    .D1(_11744_),
    .Y(_11752_));
 sky130_fd_sc_hd__o211ai_2 _21864_ (.A1(_05990_),
    .A2(_05992_),
    .B1(_11749_),
    .C1(_11752_),
    .Y(_11753_));
 sky130_fd_sc_hd__o22ai_2 _21865_ (.A1(_05990_),
    .A2(_05992_),
    .B1(_11747_),
    .B2(_11751_),
    .Y(_11754_));
 sky130_fd_sc_hd__o31a_1 _21866_ (.A1(_05990_),
    .A2(_05992_),
    .A3(_11735_),
    .B1(_11753_),
    .X(_11755_));
 sky130_fd_sc_hd__inv_2 _21867_ (.A(_11755_),
    .Y(_11756_));
 sky130_fd_sc_hd__a21oi_1 _21868_ (.A1(_11271_),
    .A2(net298),
    .B1(_11279_),
    .Y(_11757_));
 sky130_fd_sc_hd__o21ai_1 _21869_ (.A1(net298),
    .A2(_11271_),
    .B1(_11279_),
    .Y(_11758_));
 sky130_fd_sc_hd__a32oi_4 _21870_ (.A1(net299),
    .A2(_11267_),
    .A3(_11270_),
    .B1(_11278_),
    .B2(_11273_),
    .Y(_11760_));
 sky130_fd_sc_hd__a31o_1 _21871_ (.A1(net240),
    .A2(_11749_),
    .A3(_11752_),
    .B1(net294),
    .X(_11761_));
 sky130_fd_sc_hd__a311oi_1 _21872_ (.A1(net240),
    .A2(_11749_),
    .A3(_11752_),
    .B1(_11736_),
    .C1(net294),
    .Y(_11762_));
 sky130_fd_sc_hd__o211ai_2 _21873_ (.A1(net240),
    .A2(_11735_),
    .B1(net295),
    .C1(_11753_),
    .Y(_11763_));
 sky130_fd_sc_hd__a2bb2oi_2 _21874_ (.A1_N(net318),
    .A2_N(net316),
    .B1(_11738_),
    .B2(_11753_),
    .Y(_11764_));
 sky130_fd_sc_hd__o221ai_4 _21875_ (.A1(net318),
    .A2(net316),
    .B1(net240),
    .B2(_11734_),
    .C1(_11754_),
    .Y(_11765_));
 sky130_fd_sc_hd__o21a_1 _21876_ (.A1(_11736_),
    .A2(_11761_),
    .B1(_11765_),
    .X(_11766_));
 sky130_fd_sc_hd__o2111ai_1 _21877_ (.A1(net299),
    .A2(_11272_),
    .B1(_11758_),
    .C1(_11763_),
    .D1(_11765_),
    .Y(_11767_));
 sky130_fd_sc_hd__o2bb2ai_1 _21878_ (.A1_N(_11273_),
    .A2_N(_11758_),
    .B1(_11762_),
    .B2(_11764_),
    .Y(_11768_));
 sky130_fd_sc_hd__nand3_2 _21879_ (.A(_11768_),
    .B(net213),
    .C(_11767_),
    .Y(_11769_));
 sky130_fd_sc_hd__o221a_1 _21880_ (.A1(_06286_),
    .A2(_06288_),
    .B1(_11734_),
    .B2(net240),
    .C1(_11754_),
    .X(_11771_));
 sky130_fd_sc_hd__inv_2 _21881_ (.A(_11771_),
    .Y(_11772_));
 sky130_fd_sc_hd__nand3_1 _21882_ (.A(_11765_),
    .B(_11760_),
    .C(_11763_),
    .Y(_11773_));
 sky130_fd_sc_hd__o22ai_1 _21883_ (.A1(_11274_),
    .A2(_11757_),
    .B1(_11762_),
    .B2(_11764_),
    .Y(_11774_));
 sky130_fd_sc_hd__nand3_1 _21884_ (.A(_11774_),
    .B(net213),
    .C(_11773_),
    .Y(_11775_));
 sky130_fd_sc_hd__o21ai_1 _21885_ (.A1(net213),
    .A2(_11756_),
    .B1(_11769_),
    .Y(_11776_));
 sky130_fd_sc_hd__o211a_1 _21886_ (.A1(_11756_),
    .A2(net213),
    .B1(_04238_),
    .C1(_11769_),
    .X(_11777_));
 sky130_fd_sc_hd__o211ai_4 _21887_ (.A1(_11756_),
    .A2(net213),
    .B1(_04238_),
    .C1(_11769_),
    .Y(_11778_));
 sky130_fd_sc_hd__and3_1 _21888_ (.A(_11775_),
    .B(net299),
    .C(_11772_),
    .X(_11779_));
 sky130_fd_sc_hd__nand3_2 _21889_ (.A(_11775_),
    .B(net299),
    .C(_11772_),
    .Y(_11780_));
 sky130_fd_sc_hd__nand2_1 _21890_ (.A(_11778_),
    .B(_11780_),
    .Y(_11782_));
 sky130_fd_sc_hd__a22oi_1 _21891_ (.A1(_02148_),
    .A2(_11285_),
    .B1(_11295_),
    .B2(_11299_),
    .Y(_11783_));
 sky130_fd_sc_hd__o2bb2ai_2 _21892_ (.A1_N(_11295_),
    .A2_N(_11299_),
    .B1(_02137_),
    .B2(_11286_),
    .Y(_11784_));
 sky130_fd_sc_hd__o21ai_2 _21893_ (.A1(_11290_),
    .A2(_11783_),
    .B1(_11782_),
    .Y(_11785_));
 sky130_fd_sc_hd__o2111ai_4 _21894_ (.A1(_02148_),
    .A2(_11285_),
    .B1(_11778_),
    .C1(_11780_),
    .D1(_11784_),
    .Y(_11786_));
 sky130_fd_sc_hd__nand3_2 _21895_ (.A(_11785_),
    .B(_11786_),
    .C(net211),
    .Y(_11787_));
 sky130_fd_sc_hd__o211a_1 _21896_ (.A1(_11756_),
    .A2(net213),
    .B1(_06613_),
    .C1(_11769_),
    .X(_11788_));
 sky130_fd_sc_hd__or3_2 _21897_ (.A(_06608_),
    .B(net237),
    .C(_11776_),
    .X(_11789_));
 sky130_fd_sc_hd__a31o_2 _21898_ (.A1(_11785_),
    .A2(_11786_),
    .A3(net211),
    .B1(_11788_),
    .X(_11790_));
 sky130_fd_sc_hd__a22oi_4 _21899_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_11787_),
    .B2(_11789_),
    .Y(_11791_));
 sky130_fd_sc_hd__a311oi_4 _21900_ (.A1(_11785_),
    .A2(_11786_),
    .A3(net211),
    .B1(_11788_),
    .C1(_02148_),
    .Y(_11793_));
 sky130_fd_sc_hd__nand3_1 _21901_ (.A(_11787_),
    .B(_11789_),
    .C(_02137_),
    .Y(_11794_));
 sky130_fd_sc_hd__nor2_1 _21902_ (.A(_11791_),
    .B(_11793_),
    .Y(_11795_));
 sky130_fd_sc_hd__o311a_1 _21903_ (.A1(_10356_),
    .A2(_10820_),
    .A3(_10822_),
    .B1(_10825_),
    .C1(_11315_),
    .X(_11796_));
 sky130_fd_sc_hd__o22a_1 _21904_ (.A1(_11311_),
    .A2(_11305_),
    .B1(_11316_),
    .B2(_11314_),
    .X(_11797_));
 sky130_fd_sc_hd__o22ai_2 _21905_ (.A1(_11311_),
    .A2(_11305_),
    .B1(_11316_),
    .B2(_11314_),
    .Y(_11798_));
 sky130_fd_sc_hd__nand3b_1 _21906_ (.A_N(_11791_),
    .B(_11794_),
    .C(_11798_),
    .Y(_11799_));
 sky130_fd_sc_hd__o21ai_1 _21907_ (.A1(_11791_),
    .A2(_11793_),
    .B1(_11797_),
    .Y(_11800_));
 sky130_fd_sc_hd__o211ai_4 _21908_ (.A1(net230),
    .A2(_06901_),
    .B1(_11799_),
    .C1(_11800_),
    .Y(_11801_));
 sky130_fd_sc_hd__and3_1 _21909_ (.A(_06900_),
    .B(_06902_),
    .C(_11790_),
    .X(_11802_));
 sky130_fd_sc_hd__a211o_1 _21910_ (.A1(_11787_),
    .A2(_11789_),
    .B1(_06899_),
    .C1(_06901_),
    .X(_11804_));
 sky130_fd_sc_hd__o21ai_1 _21911_ (.A1(_11791_),
    .A2(_11793_),
    .B1(_11798_),
    .Y(_11805_));
 sky130_fd_sc_hd__o211a_1 _21912_ (.A1(_11314_),
    .A2(_11316_),
    .B1(_11794_),
    .C1(_11313_),
    .X(_11806_));
 sky130_fd_sc_hd__o211ai_2 _21913_ (.A1(_11314_),
    .A2(_11316_),
    .B1(_11794_),
    .C1(_11313_),
    .Y(_11807_));
 sky130_fd_sc_hd__o221ai_4 _21914_ (.A1(net230),
    .A2(_06901_),
    .B1(_11791_),
    .B2(_11807_),
    .C1(_11805_),
    .Y(_11808_));
 sky130_fd_sc_hd__o21ai_2 _21915_ (.A1(net208),
    .A2(_11790_),
    .B1(_11801_),
    .Y(_11809_));
 sky130_fd_sc_hd__inv_2 _21916_ (.A(_11809_),
    .Y(_11810_));
 sky130_fd_sc_hd__or3_2 _21917_ (.A(_07227_),
    .B(_07229_),
    .C(_11809_),
    .X(_11811_));
 sky130_fd_sc_hd__o21ai_1 _21918_ (.A1(_00218_),
    .A2(_00229_),
    .B1(_11808_),
    .Y(_11812_));
 sky130_fd_sc_hd__o211a_1 _21919_ (.A1(_00218_),
    .A2(_00229_),
    .B1(_11804_),
    .C1(_11808_),
    .X(_11813_));
 sky130_fd_sc_hd__o211ai_4 _21920_ (.A1(_00218_),
    .A2(_00229_),
    .B1(_11804_),
    .C1(_11808_),
    .Y(_11815_));
 sky130_fd_sc_hd__o211ai_4 _21921_ (.A1(_11790_),
    .A2(net208),
    .B1(_00251_),
    .C1(_11801_),
    .Y(_11816_));
 sky130_fd_sc_hd__a21oi_1 _21922_ (.A1(net326),
    .A2(_11325_),
    .B1(_11329_),
    .Y(_11817_));
 sky130_fd_sc_hd__o21ai_2 _21923_ (.A1(_11330_),
    .A2(_11333_),
    .B1(_11336_),
    .Y(_11818_));
 sky130_fd_sc_hd__a21oi_1 _21924_ (.A1(_11334_),
    .A2(_11329_),
    .B1(_11335_),
    .Y(_11819_));
 sky130_fd_sc_hd__a21oi_1 _21925_ (.A1(_11815_),
    .A2(_11816_),
    .B1(_11818_),
    .Y(_11820_));
 sky130_fd_sc_hd__o2bb2ai_2 _21926_ (.A1_N(_11815_),
    .A2_N(_11816_),
    .B1(_11817_),
    .B2(_11333_),
    .Y(_11821_));
 sky130_fd_sc_hd__o211a_1 _21927_ (.A1(_11802_),
    .A2(_11812_),
    .B1(_11816_),
    .C1(_11818_),
    .X(_11822_));
 sky130_fd_sc_hd__a31oi_4 _21928_ (.A1(_11818_),
    .A2(_11816_),
    .A3(_11815_),
    .B1(_07232_),
    .Y(_11823_));
 sky130_fd_sc_hd__nand2_2 _21929_ (.A(_11823_),
    .B(_11821_),
    .Y(_11824_));
 sky130_fd_sc_hd__o22ai_2 _21930_ (.A1(_07227_),
    .A2(_07229_),
    .B1(_11820_),
    .B2(_11822_),
    .Y(_11826_));
 sky130_fd_sc_hd__a22o_2 _21931_ (.A1(_07232_),
    .A2(_11810_),
    .B1(_11823_),
    .B2(_11821_),
    .X(_11827_));
 sky130_fd_sc_hd__a31o_1 _21932_ (.A1(_11309_),
    .A2(_11326_),
    .A3(_11339_),
    .B1(_11350_),
    .X(_11828_));
 sky130_fd_sc_hd__a22oi_2 _21933_ (.A1(_10851_),
    .A2(_10859_),
    .B1(_11345_),
    .B2(_11298_),
    .Y(_11829_));
 sky130_fd_sc_hd__a32o_1 _21934_ (.A1(_11344_),
    .A2(_11298_),
    .A3(_11340_),
    .B1(_10851_),
    .B2(_10859_),
    .X(_11830_));
 sky130_fd_sc_hd__a21o_1 _21935_ (.A1(_11348_),
    .A2(_11350_),
    .B1(_11346_),
    .X(_11831_));
 sky130_fd_sc_hd__a221oi_4 _21936_ (.A1(_07232_),
    .A2(_11810_),
    .B1(_11823_),
    .B2(_11821_),
    .C1(net326),
    .Y(_11832_));
 sky130_fd_sc_hd__o221ai_4 _21937_ (.A1(_12867_),
    .A2(_12877_),
    .B1(net185),
    .B2(_11809_),
    .C1(_11824_),
    .Y(_11833_));
 sky130_fd_sc_hd__a2bb2oi_4 _21938_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_11811_),
    .B2(_11824_),
    .Y(_11834_));
 sky130_fd_sc_hd__o211ai_4 _21939_ (.A1(_11810_),
    .A2(net185),
    .B1(net326),
    .C1(_11826_),
    .Y(_11835_));
 sky130_fd_sc_hd__nor2_1 _21940_ (.A(_11832_),
    .B(_11834_),
    .Y(_11837_));
 sky130_fd_sc_hd__o2111ai_4 _21941_ (.A1(_11298_),
    .A2(_11345_),
    .B1(_11830_),
    .C1(_11833_),
    .D1(_11835_),
    .Y(_11838_));
 sky130_fd_sc_hd__o22ai_2 _21942_ (.A1(_11346_),
    .A2(_11829_),
    .B1(_11832_),
    .B2(_11834_),
    .Y(_11839_));
 sky130_fd_sc_hd__o211ai_4 _21943_ (.A1(_07544_),
    .A2(net184),
    .B1(_11838_),
    .C1(_11839_),
    .Y(_11840_));
 sky130_fd_sc_hd__a211o_1 _21944_ (.A1(_11811_),
    .A2(_11824_),
    .B1(_07544_),
    .C1(net184),
    .X(_11841_));
 sky130_fd_sc_hd__o211ai_1 _21945_ (.A1(_11346_),
    .A2(_11829_),
    .B1(_11833_),
    .C1(_11835_),
    .Y(_11842_));
 sky130_fd_sc_hd__o2bb2ai_1 _21946_ (.A1_N(_11348_),
    .A2_N(_11828_),
    .B1(_11832_),
    .B2(_11834_),
    .Y(_11843_));
 sky130_fd_sc_hd__o211ai_2 _21947_ (.A1(_07544_),
    .A2(net184),
    .B1(_11842_),
    .C1(_11843_),
    .Y(_11844_));
 sky130_fd_sc_hd__o21ai_4 _21948_ (.A1(net163),
    .A2(_11827_),
    .B1(_11840_),
    .Y(_11845_));
 sky130_fd_sc_hd__o211a_1 _21949_ (.A1(_11827_),
    .A2(net163),
    .B1(_11309_),
    .C1(_11840_),
    .X(_11846_));
 sky130_fd_sc_hd__o211ai_4 _21950_ (.A1(_11827_),
    .A2(net163),
    .B1(_11309_),
    .C1(_11840_),
    .Y(_11848_));
 sky130_fd_sc_hd__o211ai_4 _21951_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_11841_),
    .C1(_11844_),
    .Y(_11849_));
 sky130_fd_sc_hd__inv_2 _21952_ (.A(_11849_),
    .Y(_11850_));
 sky130_fd_sc_hd__a21oi_1 _21953_ (.A1(_10025_),
    .A2(_11359_),
    .B1(_11363_),
    .Y(_11851_));
 sky130_fd_sc_hd__o21ai_1 _21954_ (.A1(_10015_),
    .A2(_11358_),
    .B1(_11371_),
    .Y(_11852_));
 sky130_fd_sc_hd__o2bb2ai_1 _21955_ (.A1_N(_11848_),
    .A2_N(_11849_),
    .B1(_11851_),
    .B2(_11367_),
    .Y(_11853_));
 sky130_fd_sc_hd__o2111ai_4 _21956_ (.A1(_11363_),
    .A2(_11365_),
    .B1(_11368_),
    .C1(_11848_),
    .D1(_11849_),
    .Y(_11854_));
 sky130_fd_sc_hd__or3_1 _21957_ (.A(_07912_),
    .B(_07914_),
    .C(_11845_),
    .X(_11855_));
 sky130_fd_sc_hd__nand3_4 _21958_ (.A(_11853_),
    .B(_11854_),
    .C(net160),
    .Y(_11856_));
 sky130_fd_sc_hd__o21ai_4 _21959_ (.A1(net160),
    .A2(_11845_),
    .B1(_11856_),
    .Y(_11857_));
 sky130_fd_sc_hd__a2bb2oi_1 _21960_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_11855_),
    .B2(_11856_),
    .Y(_11859_));
 sky130_fd_sc_hd__o21ai_4 _21961_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_11857_),
    .Y(_11860_));
 sky130_fd_sc_hd__o221a_2 _21962_ (.A1(net365),
    .A2(net362),
    .B1(net160),
    .B2(_11845_),
    .C1(_11856_),
    .X(_11861_));
 sky130_fd_sc_hd__o221ai_4 _21963_ (.A1(net365),
    .A2(net362),
    .B1(net160),
    .B2(_11845_),
    .C1(_11856_),
    .Y(_11862_));
 sky130_fd_sc_hd__a32oi_4 _21964_ (.A1(_11374_),
    .A2(_08907_),
    .A3(_11361_),
    .B1(_10885_),
    .B2(_10891_),
    .Y(_11863_));
 sky130_fd_sc_hd__a21oi_4 _21965_ (.A1(_11380_),
    .A2(_11382_),
    .B1(_11383_),
    .Y(_11864_));
 sky130_fd_sc_hd__a32o_2 _21966_ (.A1(_08874_),
    .A2(_08896_),
    .A3(_11376_),
    .B1(_11380_),
    .B2(_11382_),
    .X(_11865_));
 sky130_fd_sc_hd__o21ai_1 _21967_ (.A1(_11859_),
    .A2(_11861_),
    .B1(_11864_),
    .Y(_11866_));
 sky130_fd_sc_hd__o211ai_2 _21968_ (.A1(_11383_),
    .A2(_11863_),
    .B1(_11862_),
    .C1(_11860_),
    .Y(_11867_));
 sky130_fd_sc_hd__nand3_1 _21969_ (.A(_11860_),
    .B(_11864_),
    .C(_11862_),
    .Y(_11868_));
 sky130_fd_sc_hd__o21ai_1 _21970_ (.A1(_11859_),
    .A2(_11861_),
    .B1(_11865_),
    .Y(_11870_));
 sky130_fd_sc_hd__o211ai_2 _21971_ (.A1(net180),
    .A2(_08298_),
    .B1(_11868_),
    .C1(_11870_),
    .Y(_11871_));
 sky130_fd_sc_hd__and3_1 _21972_ (.A(_11857_),
    .B(_08299_),
    .C(_08297_),
    .X(_11872_));
 sky130_fd_sc_hd__a211o_1 _21973_ (.A1(_11855_),
    .A2(_11856_),
    .B1(net180),
    .C1(_08298_),
    .X(_11873_));
 sky130_fd_sc_hd__nand3_1 _21974_ (.A(_11866_),
    .B(_11867_),
    .C(_08300_),
    .Y(_11874_));
 sky130_fd_sc_hd__a31o_2 _21975_ (.A1(_11866_),
    .A2(_11867_),
    .A3(_08300_),
    .B1(_11872_),
    .X(_11875_));
 sky130_fd_sc_hd__a21oi_1 _21976_ (.A1(_07899_),
    .A2(_11392_),
    .B1(_11396_),
    .Y(_11876_));
 sky130_fd_sc_hd__o21ai_1 _21977_ (.A1(_11398_),
    .A2(_11399_),
    .B1(_11402_),
    .Y(_11877_));
 sky130_fd_sc_hd__a311oi_2 _21978_ (.A1(_11866_),
    .A2(_11867_),
    .A3(_08300_),
    .B1(_11872_),
    .C1(_08918_),
    .Y(_11878_));
 sky130_fd_sc_hd__o211ai_2 _21979_ (.A1(_08863_),
    .A2(_08885_),
    .B1(_11873_),
    .C1(_11874_),
    .Y(_11879_));
 sky130_fd_sc_hd__a2bb2oi_1 _21980_ (.A1_N(_08819_),
    .A2_N(_08841_),
    .B1(_11873_),
    .B2(_11874_),
    .Y(_11881_));
 sky130_fd_sc_hd__o211ai_4 _21981_ (.A1(_08300_),
    .A2(_11857_),
    .B1(_11871_),
    .C1(_08918_),
    .Y(_11882_));
 sky130_fd_sc_hd__o2111ai_1 _21982_ (.A1(_11398_),
    .A2(_11399_),
    .B1(_11402_),
    .C1(_11879_),
    .D1(_11882_),
    .Y(_11883_));
 sky130_fd_sc_hd__o22ai_1 _21983_ (.A1(_11401_),
    .A2(_11403_),
    .B1(_11878_),
    .B2(_11881_),
    .Y(_11884_));
 sky130_fd_sc_hd__nand3_2 _21984_ (.A(_11884_),
    .B(_08714_),
    .C(_11883_),
    .Y(_11885_));
 sky130_fd_sc_hd__a22o_1 _21985_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_11873_),
    .B2(_11874_),
    .X(_11886_));
 sky130_fd_sc_hd__nand3_1 _21986_ (.A(_11877_),
    .B(_11879_),
    .C(_11882_),
    .Y(_11887_));
 sky130_fd_sc_hd__o22ai_1 _21987_ (.A1(_11399_),
    .A2(_11876_),
    .B1(_11878_),
    .B2(_11881_),
    .Y(_11888_));
 sky130_fd_sc_hd__nand3_1 _21988_ (.A(_11888_),
    .B(_08714_),
    .C(_11887_),
    .Y(_11889_));
 sky130_fd_sc_hd__o21a_2 _21989_ (.A1(_08714_),
    .A2(_11875_),
    .B1(_11885_),
    .X(_11890_));
 sky130_fd_sc_hd__o211ai_4 _21990_ (.A1(_08714_),
    .A2(_11875_),
    .B1(_11885_),
    .C1(_07899_),
    .Y(_11892_));
 sky130_fd_sc_hd__nand3_4 _21991_ (.A(_11889_),
    .B(_07888_),
    .C(_11886_),
    .Y(_11893_));
 sky130_fd_sc_hd__o21a_1 _21992_ (.A1(_07033_),
    .A2(_11409_),
    .B1(_10961_),
    .X(_11894_));
 sky130_fd_sc_hd__o21ai_1 _21993_ (.A1(_07033_),
    .A2(_11409_),
    .B1(_10961_),
    .Y(_11895_));
 sky130_fd_sc_hd__o21ai_2 _21994_ (.A1(_10961_),
    .A2(_11410_),
    .B1(_11413_),
    .Y(_11896_));
 sky130_fd_sc_hd__o2bb2ai_4 _21995_ (.A1_N(_11892_),
    .A2_N(_11893_),
    .B1(_11894_),
    .B2(_11410_),
    .Y(_11897_));
 sky130_fd_sc_hd__o21ai_1 _21996_ (.A1(_07899_),
    .A2(_11890_),
    .B1(_11896_),
    .Y(_11898_));
 sky130_fd_sc_hd__a41oi_4 _21997_ (.A1(_11411_),
    .A2(_11892_),
    .A3(_11893_),
    .A4(_11895_),
    .B1(_09124_),
    .Y(_11899_));
 sky130_fd_sc_hd__o221a_2 _21998_ (.A1(_09122_),
    .A2(_09123_),
    .B1(_11875_),
    .B2(_08714_),
    .C1(_11885_),
    .X(_11900_));
 sky130_fd_sc_hd__a21oi_4 _21999_ (.A1(_11899_),
    .A2(_11897_),
    .B1(_11900_),
    .Y(_11901_));
 sky130_fd_sc_hd__a22o_1 _22000_ (.A1(_09124_),
    .A2(_11890_),
    .B1(_11899_),
    .B2(_11897_),
    .X(_11903_));
 sky130_fd_sc_hd__a21oi_2 _22001_ (.A1(_11426_),
    .A2(_11427_),
    .B1(_11424_),
    .Y(_11904_));
 sky130_fd_sc_hd__a22o_1 _22002_ (.A1(net376),
    .A2(_07022_),
    .B1(_11899_),
    .B2(_11897_),
    .X(_11905_));
 sky130_fd_sc_hd__a221oi_4 _22003_ (.A1(_09124_),
    .A2(_11890_),
    .B1(_11899_),
    .B2(_11897_),
    .C1(_07044_),
    .Y(_11906_));
 sky130_fd_sc_hd__a21oi_2 _22004_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_11901_),
    .Y(_11907_));
 sky130_fd_sc_hd__o21ai_4 _22005_ (.A1(_06945_),
    .A2(_06967_),
    .B1(_11903_),
    .Y(_11908_));
 sky130_fd_sc_hd__o221ai_4 _22006_ (.A1(_11900_),
    .A2(_11905_),
    .B1(_11424_),
    .B2(_11429_),
    .C1(_11908_),
    .Y(_11909_));
 sky130_fd_sc_hd__o21ai_1 _22007_ (.A1(_11906_),
    .A2(_11907_),
    .B1(_11904_),
    .Y(_11910_));
 sky130_fd_sc_hd__or3_1 _22008_ (.A(_09553_),
    .B(net155),
    .C(_11901_),
    .X(_11911_));
 sky130_fd_sc_hd__o2111ai_4 _22009_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .C1(_11909_),
    .D1(_11910_),
    .Y(_11912_));
 sky130_fd_sc_hd__a21oi_2 _22010_ (.A1(_11911_),
    .A2(_11912_),
    .B1(_06332_),
    .Y(_11914_));
 sky130_fd_sc_hd__o221a_1 _22011_ (.A1(net381),
    .A2(_06310_),
    .B1(net143),
    .B2(_11901_),
    .C1(_11912_),
    .X(_11915_));
 sky130_fd_sc_hd__o221ai_4 _22012_ (.A1(net381),
    .A2(_06310_),
    .B1(net143),
    .B2(_11901_),
    .C1(_11912_),
    .Y(_11916_));
 sky130_fd_sc_hd__a31oi_2 _22013_ (.A1(_11423_),
    .A2(_11432_),
    .A3(_11435_),
    .B1(_11436_),
    .Y(_11917_));
 sky130_fd_sc_hd__o21bai_1 _22014_ (.A1(_11914_),
    .A2(_11915_),
    .B1_N(_11917_),
    .Y(_11918_));
 sky130_fd_sc_hd__nand2_1 _22015_ (.A(_11916_),
    .B(_11917_),
    .Y(_11919_));
 sky130_fd_sc_hd__o21ai_1 _22016_ (.A1(_11914_),
    .A2(_11919_),
    .B1(_11918_),
    .Y(_11920_));
 sky130_fd_sc_hd__o311a_1 _22017_ (.A1(_09553_),
    .A2(net155),
    .A3(_11901_),
    .B1(_09578_),
    .C1(_11912_),
    .X(_11921_));
 sky130_fd_sc_hd__a21oi_2 _22018_ (.A1(_11920_),
    .A2(_09579_),
    .B1(_11921_),
    .Y(_11922_));
 sky130_fd_sc_hd__a32oi_4 _22019_ (.A1(_05512_),
    .A2(net396),
    .A3(_11442_),
    .B1(_11440_),
    .B2(_11444_),
    .Y(_11923_));
 sky130_fd_sc_hd__and3_1 _22020_ (.A(_11923_),
    .B(_05796_),
    .C(net395),
    .X(_11925_));
 sky130_fd_sc_hd__a21oi_1 _22021_ (.A1(net395),
    .A2(_05796_),
    .B1(_11923_),
    .Y(_11926_));
 sky130_fd_sc_hd__o21ai_2 _22022_ (.A1(_05851_),
    .A2(_11923_),
    .B1(_10480_),
    .Y(_11927_));
 sky130_fd_sc_hd__o21ai_1 _22023_ (.A1(_11927_),
    .A2(_11925_),
    .B1(_11922_),
    .Y(_11928_));
 sky130_fd_sc_hd__o31ai_4 _22024_ (.A1(_11925_),
    .A2(_11927_),
    .A3(_11922_),
    .B1(_11928_),
    .Y(_11929_));
 sky130_fd_sc_hd__a211o_1 _22025_ (.A1(_05512_),
    .A2(net396),
    .B1(_11448_),
    .C1(_11450_),
    .X(_11930_));
 sky130_fd_sc_hd__o221a_1 _22026_ (.A1(_03399_),
    .A2(_05491_),
    .B1(_11448_),
    .B2(_11450_),
    .C1(net396),
    .X(_11931_));
 sky130_fd_sc_hd__o21ai_1 _22027_ (.A1(_11448_),
    .A2(_11450_),
    .B1(_05556_),
    .Y(_11932_));
 sky130_fd_sc_hd__nand2_1 _22028_ (.A(_11930_),
    .B(_11932_),
    .Y(_11933_));
 sky130_fd_sc_hd__o21ai_1 _22029_ (.A1(_10953_),
    .A2(_11933_),
    .B1(_11929_),
    .Y(_11934_));
 sky130_fd_sc_hd__o31a_1 _22030_ (.A1(_10953_),
    .A2(_11929_),
    .A3(_11933_),
    .B1(_11934_),
    .X(_11936_));
 sky130_fd_sc_hd__or3_1 _22031_ (.A(net407),
    .B(_05218_),
    .C(_11936_),
    .X(_11937_));
 sky130_fd_sc_hd__o311ai_2 _22032_ (.A1(_10953_),
    .A2(_11929_),
    .A3(_11933_),
    .B1(_11934_),
    .C1(_05250_),
    .Y(_11938_));
 sky130_fd_sc_hd__nand2_1 _22033_ (.A(_11937_),
    .B(_11938_),
    .Y(_11939_));
 sky130_fd_sc_hd__nand2_1 _22034_ (.A(_11456_),
    .B(_11938_),
    .Y(_11940_));
 sky130_fd_sc_hd__xor2_1 _22035_ (.A(_11456_),
    .B(_11939_),
    .X(_11941_));
 sky130_fd_sc_hd__mux2_1 _22036_ (.A0(_11941_),
    .A1(_11936_),
    .S(_11464_),
    .X(_11942_));
 sky130_fd_sc_hd__nor4b_4 _22037_ (.A(net54),
    .B(net56),
    .C(_10947_),
    .D_N(net57),
    .Y(_11943_));
 sky130_fd_sc_hd__or4b_4 _22038_ (.A(net54),
    .B(net56),
    .C(_10947_),
    .D_N(net57),
    .X(_11944_));
 sky130_fd_sc_hd__o21ai_2 _22039_ (.A1(_03289_),
    .A2(_11944_),
    .B1(_11942_),
    .Y(_11945_));
 sky130_fd_sc_hd__and3_1 _22040_ (.A(_05119_),
    .B(_11468_),
    .C(_11945_),
    .X(_11947_));
 sky130_fd_sc_hd__a21oi_1 _22041_ (.A1(_05119_),
    .A2(_11468_),
    .B1(_11945_),
    .Y(_11948_));
 sky130_fd_sc_hd__nor2_1 _22042_ (.A(_11947_),
    .B(_11948_),
    .Y(net89));
 sky130_fd_sc_hd__o22a_1 _22043_ (.A1(_04832_),
    .A2(_04942_),
    .B1(_11468_),
    .B2(_11945_),
    .X(_11949_));
 sky130_fd_sc_hd__o21ai_1 _22044_ (.A1(_08918_),
    .A2(_11875_),
    .B1(_11877_),
    .Y(_11950_));
 sky130_fd_sc_hd__a21o_2 _22045_ (.A1(_11877_),
    .A2(_11879_),
    .B1(_11881_),
    .X(_11951_));
 sky130_fd_sc_hd__nand4_2 _22046_ (.A(_10368_),
    .B(_10370_),
    .C(_10840_),
    .D(_10842_),
    .Y(_11952_));
 sky130_fd_sc_hd__a21oi_1 _22047_ (.A1(net326),
    .A2(_11325_),
    .B1(_11952_),
    .Y(_11953_));
 sky130_fd_sc_hd__a211oi_2 _22048_ (.A1(_11332_),
    .A2(_11310_),
    .B1(_11952_),
    .C1(_11335_),
    .Y(_11954_));
 sky130_fd_sc_hd__nand3_1 _22049_ (.A(_11953_),
    .B(_11815_),
    .C(_11334_),
    .Y(_11955_));
 sky130_fd_sc_hd__o211ai_4 _22050_ (.A1(_11819_),
    .A2(_11813_),
    .B1(_11816_),
    .C1(_11955_),
    .Y(_11957_));
 sky130_fd_sc_hd__nand4b_4 _22051_ (.A_N(_10371_),
    .B(_11954_),
    .C(_11816_),
    .D(_11815_),
    .Y(_11958_));
 sky130_fd_sc_hd__nand2_1 _22052_ (.A(_11957_),
    .B(_11958_),
    .Y(_11959_));
 sky130_fd_sc_hd__o21a_1 _22053_ (.A1(_05185_),
    .A2(_11471_),
    .B1(_10970_),
    .X(_11960_));
 sky130_fd_sc_hd__and3_1 _22054_ (.A(_11476_),
    .B(_05163_),
    .C(_05141_),
    .X(_11961_));
 sky130_fd_sc_hd__a31o_1 _22055_ (.A1(_11476_),
    .A2(_05163_),
    .A3(_05141_),
    .B1(_11960_),
    .X(_11962_));
 sky130_fd_sc_hd__a21boi_1 _22056_ (.A1(_11485_),
    .A2(_11482_),
    .B1_N(_11480_),
    .Y(_11963_));
 sky130_fd_sc_hd__o211ai_2 _22057_ (.A1(_11960_),
    .A2(_11961_),
    .B1(_11480_),
    .C1(_11486_),
    .Y(_11964_));
 sky130_fd_sc_hd__a21oi_1 _22058_ (.A1(_11480_),
    .A2(_11486_),
    .B1(_11962_),
    .Y(_11965_));
 sky130_fd_sc_hd__o2111ai_4 _22059_ (.A1(_11470_),
    .A2(_11476_),
    .B1(net405),
    .C1(_05359_),
    .D1(_05381_),
    .Y(_11966_));
 sky130_fd_sc_hd__o221ai_4 _22060_ (.A1(_05348_),
    .A2(net401),
    .B1(_11962_),
    .B2(_11963_),
    .C1(_11964_),
    .Y(_11968_));
 sky130_fd_sc_hd__and2_1 _22061_ (.A(_11966_),
    .B(_11968_),
    .X(_11969_));
 sky130_fd_sc_hd__or3_1 _22062_ (.A(_05676_),
    .B(_05698_),
    .C(_11969_),
    .X(_11970_));
 sky130_fd_sc_hd__inv_2 _22063_ (.A(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__a2bb2oi_1 _22064_ (.A1_N(_10487_),
    .A2_N(_10488_),
    .B1(_11966_),
    .B2(_11968_),
    .Y(_11972_));
 sky130_fd_sc_hd__a2bb2o_1 _22065_ (.A1_N(_10487_),
    .A2_N(_10488_),
    .B1(_11966_),
    .B2(_11968_),
    .X(_11973_));
 sky130_fd_sc_hd__o211a_1 _22066_ (.A1(_10489_),
    .A2(_10490_),
    .B1(_11966_),
    .C1(_11968_),
    .X(_11974_));
 sky130_fd_sc_hd__o211ai_1 _22067_ (.A1(_10489_),
    .A2(_10490_),
    .B1(_11966_),
    .C1(_11968_),
    .Y(_11975_));
 sky130_fd_sc_hd__nand2_2 _22068_ (.A(_11973_),
    .B(_11975_),
    .Y(_11976_));
 sky130_fd_sc_hd__o32a_1 _22069_ (.A1(_11508_),
    .A2(_11499_),
    .A3(_11505_),
    .B1(_11490_),
    .B2(_10026_),
    .X(_11977_));
 sky130_fd_sc_hd__a21oi_4 _22070_ (.A1(_11494_),
    .A2(_11513_),
    .B1(_11976_),
    .Y(_11979_));
 sky130_fd_sc_hd__o22ai_2 _22071_ (.A1(_10026_),
    .A2(_11490_),
    .B1(_11972_),
    .B2(_11974_),
    .Y(_11980_));
 sky130_fd_sc_hd__o22ai_4 _22072_ (.A1(_05676_),
    .A2(_05698_),
    .B1(_11980_),
    .B2(_11512_),
    .Y(_11981_));
 sky130_fd_sc_hd__o22a_2 _22073_ (.A1(net358),
    .A2(_11969_),
    .B1(_11981_),
    .B2(_11979_),
    .X(_11982_));
 sky130_fd_sc_hd__o22ai_4 _22074_ (.A1(net358),
    .A2(_11969_),
    .B1(_11981_),
    .B2(_11979_),
    .Y(_11983_));
 sky130_fd_sc_hd__and3_1 _22075_ (.A(_06804_),
    .B(_06826_),
    .C(_11983_),
    .X(_11984_));
 sky130_fd_sc_hd__or3_2 _22076_ (.A(_06793_),
    .B(_06815_),
    .C(_11982_),
    .X(_11985_));
 sky130_fd_sc_hd__o21a_1 _22077_ (.A1(_10021_),
    .A2(_10022_),
    .B1(_11983_),
    .X(_11986_));
 sky130_fd_sc_hd__o21ai_2 _22078_ (.A1(_10021_),
    .A2(_10022_),
    .B1(_11983_),
    .Y(_11987_));
 sky130_fd_sc_hd__o21ai_2 _22079_ (.A1(_11981_),
    .A2(_11979_),
    .B1(_10026_),
    .Y(_11988_));
 sky130_fd_sc_hd__o221a_1 _22080_ (.A1(net358),
    .A2(_11969_),
    .B1(_11981_),
    .B2(_11979_),
    .C1(_10026_),
    .X(_11990_));
 sky130_fd_sc_hd__o21a_2 _22081_ (.A1(_11971_),
    .A2(_11988_),
    .B1(_11987_),
    .X(_11991_));
 sky130_fd_sc_hd__o21ai_4 _22082_ (.A1(_11971_),
    .A2(_11988_),
    .B1(_11987_),
    .Y(_11992_));
 sky130_fd_sc_hd__nand3_1 _22083_ (.A(_10543_),
    .B(_10545_),
    .C(_10081_),
    .Y(_11993_));
 sky130_fd_sc_hd__nor3_1 _22084_ (.A(_11028_),
    .B(_11030_),
    .C(_11993_),
    .Y(_11994_));
 sky130_fd_sc_hd__a21oi_4 _22085_ (.A1(_11994_),
    .A2(_11524_),
    .B1(_11520_),
    .Y(_11995_));
 sky130_fd_sc_hd__nand2_1 _22086_ (.A(_11529_),
    .B(_11995_),
    .Y(_11996_));
 sky130_fd_sc_hd__and4b_1 _22087_ (.A_N(_11993_),
    .B(_11031_),
    .C(_11029_),
    .D(_10093_),
    .X(_11997_));
 sky130_fd_sc_hd__nand4b_4 _22088_ (.A_N(_11993_),
    .B(_11031_),
    .C(_11029_),
    .D(_10093_),
    .Y(_11998_));
 sky130_fd_sc_hd__nor3_1 _22089_ (.A(_11998_),
    .B(_11523_),
    .C(_11520_),
    .Y(_11999_));
 sky130_fd_sc_hd__a22oi_4 _22090_ (.A1(_11525_),
    .A2(_11997_),
    .B1(_11529_),
    .B2(_11995_),
    .Y(_12001_));
 sky130_fd_sc_hd__o2bb2ai_4 _22091_ (.A1_N(_11995_),
    .A2_N(_11529_),
    .B1(_11526_),
    .B2(_11998_),
    .Y(_12002_));
 sky130_fd_sc_hd__o21ai_2 _22092_ (.A1(_11986_),
    .A2(_11990_),
    .B1(_12002_),
    .Y(_12003_));
 sky130_fd_sc_hd__a211oi_4 _22093_ (.A1(_11529_),
    .A2(_11995_),
    .B1(_11999_),
    .C1(_11992_),
    .Y(_12004_));
 sky130_fd_sc_hd__o211ai_2 _22094_ (.A1(_11526_),
    .A2(_11998_),
    .B1(_11991_),
    .C1(_11996_),
    .Y(_12005_));
 sky130_fd_sc_hd__o22ai_4 _22095_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_11991_),
    .B2(_12001_),
    .Y(_12006_));
 sky130_fd_sc_hd__o221ai_4 _22096_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_11992_),
    .B2(_12002_),
    .C1(_12003_),
    .Y(_12007_));
 sky130_fd_sc_hd__o22ai_1 _22097_ (.A1(net357),
    .A2(_11982_),
    .B1(_12004_),
    .B2(_12006_),
    .Y(_12008_));
 sky130_fd_sc_hd__a21oi_2 _22098_ (.A1(_11985_),
    .A2(_12007_),
    .B1(net354),
    .Y(_12009_));
 sky130_fd_sc_hd__a211o_1 _22099_ (.A1(_11985_),
    .A2(_12007_),
    .B1(net374),
    .C1(_07702_),
    .X(_12010_));
 sky130_fd_sc_hd__o221ai_4 _22100_ (.A1(net174),
    .A2(_11532_),
    .B1(_11047_),
    .B2(_11048_),
    .C1(_11043_),
    .Y(_12012_));
 sky130_fd_sc_hd__a311oi_4 _22101_ (.A1(_12003_),
    .A2(_12005_),
    .A3(net357),
    .B1(_09595_),
    .C1(_11984_),
    .Y(_12013_));
 sky130_fd_sc_hd__o221ai_4 _22102_ (.A1(net357),
    .A2(_11982_),
    .B1(_12004_),
    .B2(_12006_),
    .C1(net172),
    .Y(_12014_));
 sky130_fd_sc_hd__a2bb2oi_4 _22103_ (.A1_N(_09588_),
    .A2_N(net187),
    .B1(_11985_),
    .B2(_12007_),
    .Y(_12015_));
 sky130_fd_sc_hd__o21ai_1 _22104_ (.A1(_09588_),
    .A2(net187),
    .B1(_12008_),
    .Y(_12016_));
 sky130_fd_sc_hd__nand4_4 _22105_ (.A(_11535_),
    .B(_12012_),
    .C(_12014_),
    .D(_12016_),
    .Y(_12017_));
 sky130_fd_sc_hd__o2bb2ai_4 _22106_ (.A1_N(_11535_),
    .A2_N(_12012_),
    .B1(_12013_),
    .B2(_12015_),
    .Y(_12018_));
 sky130_fd_sc_hd__nand3_1 _22107_ (.A(_12017_),
    .B(_12018_),
    .C(net354),
    .Y(_12019_));
 sky130_fd_sc_hd__a31oi_4 _22108_ (.A1(_12017_),
    .A2(_12018_),
    .A3(net354),
    .B1(_12009_),
    .Y(_12020_));
 sky130_fd_sc_hd__a31o_2 _22109_ (.A1(_12017_),
    .A2(_12018_),
    .A3(net354),
    .B1(_12009_),
    .X(_12021_));
 sky130_fd_sc_hd__a2bb2oi_2 _22110_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_12010_),
    .B2(_12019_),
    .Y(_12023_));
 sky130_fd_sc_hd__a2bb2o_1 _22111_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_12010_),
    .B2(_12019_),
    .X(_12024_));
 sky130_fd_sc_hd__a31oi_1 _22112_ (.A1(_12017_),
    .A2(_12018_),
    .A3(net354),
    .B1(net173),
    .Y(_12025_));
 sky130_fd_sc_hd__and3_2 _22113_ (.A(_12019_),
    .B(net174),
    .C(_12010_),
    .X(_12026_));
 sky130_fd_sc_hd__a311o_1 _22114_ (.A1(_12017_),
    .A2(_12018_),
    .A3(net354),
    .B1(net173),
    .C1(_12009_),
    .X(_12027_));
 sky130_fd_sc_hd__a21oi_1 _22115_ (.A1(_12010_),
    .A2(_12025_),
    .B1(_12023_),
    .Y(_12028_));
 sky130_fd_sc_hd__nand2_1 _22116_ (.A(_12024_),
    .B(_12027_),
    .Y(_12029_));
 sky130_fd_sc_hd__o31ai_1 _22117_ (.A1(_11056_),
    .A2(_11548_),
    .A3(_11551_),
    .B1(_11547_),
    .Y(_12030_));
 sky130_fd_sc_hd__o221a_1 _22118_ (.A1(_11548_),
    .A2(_11554_),
    .B1(_12023_),
    .B2(_12026_),
    .C1(_11547_),
    .X(_12031_));
 sky130_fd_sc_hd__o221ai_2 _22119_ (.A1(_11548_),
    .A2(_11554_),
    .B1(_12023_),
    .B2(_12026_),
    .C1(_11547_),
    .Y(_12032_));
 sky130_fd_sc_hd__a21oi_1 _22120_ (.A1(_11547_),
    .A2(_11555_),
    .B1(_12029_),
    .Y(_12034_));
 sky130_fd_sc_hd__nand2_1 _22121_ (.A(_12030_),
    .B(_12028_),
    .Y(_12035_));
 sky130_fd_sc_hd__o22ai_2 _22122_ (.A1(_08678_),
    .A2(_08700_),
    .B1(_12031_),
    .B2(_12034_),
    .Y(_12036_));
 sky130_fd_sc_hd__or3_1 _22123_ (.A(_08678_),
    .B(_08700_),
    .C(_12020_),
    .X(_12037_));
 sky130_fd_sc_hd__nand3_2 _22124_ (.A(_12035_),
    .B(net338),
    .C(_12032_),
    .Y(_12038_));
 sky130_fd_sc_hd__o31a_2 _22125_ (.A1(_08678_),
    .A2(_08700_),
    .A3(_12020_),
    .B1(_12038_),
    .X(_12039_));
 sky130_fd_sc_hd__or3_2 _22126_ (.A(net351),
    .B(_09807_),
    .C(_12039_),
    .X(_12040_));
 sky130_fd_sc_hd__a2bb2oi_2 _22127_ (.A1_N(_08724_),
    .A2_N(_08726_),
    .B1(_12037_),
    .B2(_12038_),
    .Y(_12041_));
 sky130_fd_sc_hd__o221ai_4 _22128_ (.A1(_08724_),
    .A2(_08726_),
    .B1(_12021_),
    .B2(net338),
    .C1(_12036_),
    .Y(_12042_));
 sky130_fd_sc_hd__o211a_2 _22129_ (.A1(net338),
    .A2(_12020_),
    .B1(net177),
    .C1(_12038_),
    .X(_12043_));
 sky130_fd_sc_hd__o211ai_4 _22130_ (.A1(net338),
    .A2(_12020_),
    .B1(net177),
    .C1(_12038_),
    .Y(_12045_));
 sky130_fd_sc_hd__a2bb2oi_1 _22131_ (.A1_N(net199),
    .A2_N(_11560_),
    .B1(_11575_),
    .B2(_11577_),
    .Y(_12046_));
 sky130_fd_sc_hd__o41ai_2 _22132_ (.A1(_08311_),
    .A2(_08312_),
    .A3(_11558_),
    .A4(_11559_),
    .B1(_11579_),
    .Y(_12047_));
 sky130_fd_sc_hd__a31oi_2 _22133_ (.A1(_11567_),
    .A2(_11575_),
    .A3(_11577_),
    .B1(_11563_),
    .Y(_12048_));
 sky130_fd_sc_hd__o2111ai_4 _22134_ (.A1(net198),
    .A2(_11562_),
    .B1(_12042_),
    .C1(_12045_),
    .D1(_12047_),
    .Y(_12049_));
 sky130_fd_sc_hd__o211ai_4 _22135_ (.A1(_12041_),
    .A2(_12043_),
    .B1(_11564_),
    .C1(_11582_),
    .Y(_12050_));
 sky130_fd_sc_hd__nand3_4 _22136_ (.A(_12049_),
    .B(_12050_),
    .C(net335),
    .Y(_12051_));
 sky130_fd_sc_hd__o31a_1 _22137_ (.A1(net351),
    .A2(_09807_),
    .A3(_12039_),
    .B1(_12051_),
    .X(_12052_));
 sky130_fd_sc_hd__inv_2 _22138_ (.A(_12052_),
    .Y(_12053_));
 sky130_fd_sc_hd__and3_1 _22139_ (.A(_10155_),
    .B(_10615_),
    .C(_10616_),
    .X(_12054_));
 sky130_fd_sc_hd__nand3_1 _22140_ (.A(_11596_),
    .B(_12054_),
    .C(_11107_),
    .Y(_12056_));
 sky130_fd_sc_hd__o211ai_4 _22141_ (.A1(_11593_),
    .A2(_11595_),
    .B1(_11598_),
    .C1(_12056_),
    .Y(_12057_));
 sky130_fd_sc_hd__and4_1 _22142_ (.A(_11103_),
    .B(_12054_),
    .C(_11106_),
    .D(_10165_),
    .X(_12058_));
 sky130_fd_sc_hd__nand3_4 _22143_ (.A(_12058_),
    .B(_11598_),
    .C(_11596_),
    .Y(_12059_));
 sky130_fd_sc_hd__nand2_4 _22144_ (.A(_12057_),
    .B(_12059_),
    .Y(_12060_));
 sky130_fd_sc_hd__a2bb2oi_4 _22145_ (.A1_N(_08307_),
    .A2_N(_08309_),
    .B1(_12040_),
    .B2(_12051_),
    .Y(_12061_));
 sky130_fd_sc_hd__a22o_2 _22146_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_12040_),
    .B2(_12051_),
    .X(_12062_));
 sky130_fd_sc_hd__a31oi_2 _22147_ (.A1(_12049_),
    .A2(_12050_),
    .A3(net335),
    .B1(net198),
    .Y(_12063_));
 sky130_fd_sc_hd__o221a_2 _22148_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_12039_),
    .B2(net335),
    .C1(_12051_),
    .X(_12064_));
 sky130_fd_sc_hd__o21ai_4 _22149_ (.A1(net335),
    .A2(_12039_),
    .B1(_12063_),
    .Y(_12065_));
 sky130_fd_sc_hd__a21oi_1 _22150_ (.A1(_12040_),
    .A2(_12063_),
    .B1(_12061_),
    .Y(_12067_));
 sky130_fd_sc_hd__nand2_1 _22151_ (.A(_12060_),
    .B(_12067_),
    .Y(_12068_));
 sky130_fd_sc_hd__o211ai_1 _22152_ (.A1(_12061_),
    .A2(_12064_),
    .B1(_12057_),
    .C1(_12059_),
    .Y(_12069_));
 sky130_fd_sc_hd__o2bb2ai_2 _22153_ (.A1_N(_12057_),
    .A2_N(_12059_),
    .B1(_12061_),
    .B2(_12064_),
    .Y(_12070_));
 sky130_fd_sc_hd__nand4_4 _22154_ (.A(_12057_),
    .B(_12059_),
    .C(_12062_),
    .D(_12065_),
    .Y(_12071_));
 sky130_fd_sc_hd__nand3_2 _22155_ (.A(_12068_),
    .B(_12069_),
    .C(net332),
    .Y(_12072_));
 sky130_fd_sc_hd__a21oi_2 _22156_ (.A1(_12040_),
    .A2(_12051_),
    .B1(net332),
    .Y(_12073_));
 sky130_fd_sc_hd__or3_1 _22157_ (.A(_11046_),
    .B(_11057_),
    .C(_12052_),
    .X(_12074_));
 sky130_fd_sc_hd__nand3_1 _22158_ (.A(_12070_),
    .B(_12071_),
    .C(net332),
    .Y(_12075_));
 sky130_fd_sc_hd__a31o_1 _22159_ (.A1(_12070_),
    .A2(_12071_),
    .A3(net332),
    .B1(_12073_),
    .X(_12076_));
 sky130_fd_sc_hd__a31oi_2 _22160_ (.A1(_12070_),
    .A2(_12071_),
    .A3(net332),
    .B1(_12073_),
    .Y(_12078_));
 sky130_fd_sc_hd__o211a_1 _22161_ (.A1(_12053_),
    .A2(net332),
    .B1(_12703_),
    .C1(_12072_),
    .X(_12079_));
 sky130_fd_sc_hd__or3_1 _22162_ (.A(net329),
    .B(net327),
    .C(_12078_),
    .X(_12080_));
 sky130_fd_sc_hd__o211ai_4 _22163_ (.A1(_12053_),
    .A2(net332),
    .B1(_07936_),
    .C1(_12072_),
    .Y(_12081_));
 sky130_fd_sc_hd__a311oi_4 _22164_ (.A1(_12070_),
    .A2(_12071_),
    .A3(net332),
    .B1(_12073_),
    .C1(_07936_),
    .Y(_12082_));
 sky130_fd_sc_hd__nand3_4 _22165_ (.A(_12075_),
    .B(_07935_),
    .C(_12074_),
    .Y(_12083_));
 sky130_fd_sc_hd__o211a_1 _22166_ (.A1(_11118_),
    .A2(net222),
    .B1(_11613_),
    .C1(_11609_),
    .X(_12084_));
 sky130_fd_sc_hd__o211ai_1 _22167_ (.A1(_11118_),
    .A2(net222),
    .B1(_11613_),
    .C1(_11609_),
    .Y(_12085_));
 sky130_fd_sc_hd__a31o_1 _22168_ (.A1(_11122_),
    .A2(_11609_),
    .A3(_11613_),
    .B1(_11610_),
    .X(_12086_));
 sky130_fd_sc_hd__a31oi_2 _22169_ (.A1(_11122_),
    .A2(_11609_),
    .A3(_11613_),
    .B1(_11610_),
    .Y(_12087_));
 sky130_fd_sc_hd__a21oi_2 _22170_ (.A1(_12081_),
    .A2(_12083_),
    .B1(_12086_),
    .Y(_12089_));
 sky130_fd_sc_hd__a21o_1 _22171_ (.A1(_12081_),
    .A2(_12083_),
    .B1(_12086_),
    .X(_12090_));
 sky130_fd_sc_hd__o2bb2ai_1 _22172_ (.A1_N(_11611_),
    .A2_N(_12085_),
    .B1(_07935_),
    .B2(_12078_),
    .Y(_12091_));
 sky130_fd_sc_hd__o211a_1 _22173_ (.A1(_11610_),
    .A2(_12084_),
    .B1(_12083_),
    .C1(_12081_),
    .X(_12092_));
 sky130_fd_sc_hd__o22ai_2 _22174_ (.A1(net329),
    .A2(net327),
    .B1(_12082_),
    .B2(_12091_),
    .Y(_12093_));
 sky130_fd_sc_hd__o211ai_1 _22175_ (.A1(_12082_),
    .A2(_12091_),
    .B1(net311),
    .C1(_12090_),
    .Y(_12094_));
 sky130_fd_sc_hd__o22ai_2 _22176_ (.A1(net329),
    .A2(net327),
    .B1(_12089_),
    .B2(_12092_),
    .Y(_12095_));
 sky130_fd_sc_hd__o22a_1 _22177_ (.A1(net311),
    .A2(_12078_),
    .B1(_12089_),
    .B2(_12093_),
    .X(_12096_));
 sky130_fd_sc_hd__a22oi_2 _22178_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_12080_),
    .B2(_12094_),
    .Y(_12097_));
 sky130_fd_sc_hd__o221ai_4 _22179_ (.A1(_07555_),
    .A2(net218),
    .B1(_12076_),
    .B2(net311),
    .C1(_12095_),
    .Y(_12098_));
 sky130_fd_sc_hd__o22ai_2 _22180_ (.A1(_07560_),
    .A2(_07562_),
    .B1(_12089_),
    .B2(_12093_),
    .Y(_12100_));
 sky130_fd_sc_hd__o221a_2 _22181_ (.A1(net311),
    .A2(_12078_),
    .B1(_12089_),
    .B2(_12093_),
    .C1(_07564_),
    .X(_12101_));
 sky130_fd_sc_hd__o22ai_1 _22182_ (.A1(net224),
    .A2(_11624_),
    .B1(_11630_),
    .B2(_11632_),
    .Y(_12102_));
 sky130_fd_sc_hd__o221ai_4 _22183_ (.A1(_11624_),
    .A2(net224),
    .B1(_12101_),
    .B2(_12097_),
    .C1(_11634_),
    .Y(_12103_));
 sky130_fd_sc_hd__o211ai_2 _22184_ (.A1(_12100_),
    .A2(_12079_),
    .B1(_12098_),
    .C1(_12102_),
    .Y(_12104_));
 sky130_fd_sc_hd__or3_1 _22185_ (.A(_00011_),
    .B(net323),
    .C(_12096_),
    .X(_12105_));
 sky130_fd_sc_hd__nand3_4 _22186_ (.A(_12103_),
    .B(_12104_),
    .C(net308),
    .Y(_12106_));
 sky130_fd_sc_hd__a2bb2oi_1 _22187_ (.A1_N(_07242_),
    .A2_N(_07243_),
    .B1(_12105_),
    .B2(_12106_),
    .Y(_12107_));
 sky130_fd_sc_hd__a2bb2o_2 _22188_ (.A1_N(_07242_),
    .A2_N(_07243_),
    .B1(_12105_),
    .B2(_12106_),
    .X(_12108_));
 sky130_fd_sc_hd__o211a_2 _22189_ (.A1(net307),
    .A2(_12096_),
    .B1(net224),
    .C1(_12106_),
    .X(_12109_));
 sky130_fd_sc_hd__o211ai_2 _22190_ (.A1(net307),
    .A2(_12096_),
    .B1(net224),
    .C1(_12106_),
    .Y(_12111_));
 sky130_fd_sc_hd__a32oi_4 _22191_ (.A1(_11655_),
    .A2(_11164_),
    .A3(_11162_),
    .B1(net227),
    .B2(_11637_),
    .Y(_12112_));
 sky130_fd_sc_hd__o21ai_1 _22192_ (.A1(net225),
    .A2(_11639_),
    .B1(_11657_),
    .Y(_12113_));
 sky130_fd_sc_hd__o22ai_1 _22193_ (.A1(net227),
    .A2(_11637_),
    .B1(_12113_),
    .B2(_11653_),
    .Y(_12114_));
 sky130_fd_sc_hd__a22oi_4 _22194_ (.A1(net225),
    .A2(_11639_),
    .B1(_12112_),
    .B2(_11654_),
    .Y(_12115_));
 sky130_fd_sc_hd__nand3_2 _22195_ (.A(_12114_),
    .B(_12111_),
    .C(_12108_),
    .Y(_12116_));
 sky130_fd_sc_hd__o21ai_2 _22196_ (.A1(_12107_),
    .A2(_12109_),
    .B1(_12115_),
    .Y(_12117_));
 sky130_fd_sc_hd__a211o_4 _22197_ (.A1(_12105_),
    .A2(_12106_),
    .B1(net304),
    .C1(_01951_),
    .X(_12118_));
 sky130_fd_sc_hd__nand3_4 _22198_ (.A(_12116_),
    .B(_12117_),
    .C(net279),
    .Y(_12119_));
 sky130_fd_sc_hd__and2_1 _22199_ (.A(_12118_),
    .B(_12119_),
    .X(_12120_));
 sky130_fd_sc_hd__a21oi_4 _22200_ (.A1(_12118_),
    .A2(_12119_),
    .B1(net277),
    .Y(_12122_));
 sky130_fd_sc_hd__a211o_1 _22201_ (.A1(_12118_),
    .A2(_12119_),
    .B1(net302),
    .C1(_04019_),
    .X(_12123_));
 sky130_fd_sc_hd__a2bb2oi_4 _22202_ (.A1_N(_06914_),
    .A2_N(_06916_),
    .B1(_12118_),
    .B2(_12119_),
    .Y(_12124_));
 sky130_fd_sc_hd__a22o_2 _22203_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_12118_),
    .B2(_12119_),
    .X(_12125_));
 sky130_fd_sc_hd__a31oi_2 _22204_ (.A1(_12116_),
    .A2(_12117_),
    .A3(net279),
    .B1(net225),
    .Y(_12126_));
 sky130_fd_sc_hd__and3_1 _22205_ (.A(_12119_),
    .B(net227),
    .C(_12118_),
    .X(_12127_));
 sky130_fd_sc_hd__nand2_2 _22206_ (.A(_12126_),
    .B(_12118_),
    .Y(_12128_));
 sky130_fd_sc_hd__a21oi_2 _22207_ (.A1(_12118_),
    .A2(_12126_),
    .B1(_12124_),
    .Y(_12129_));
 sky130_fd_sc_hd__nand4_2 _22208_ (.A(_10219_),
    .B(_10220_),
    .C(_10691_),
    .D(_10693_),
    .Y(_12130_));
 sky130_fd_sc_hd__a211oi_4 _22209_ (.A1(_11160_),
    .A2(_11176_),
    .B1(_12130_),
    .C1(_11180_),
    .Y(_12131_));
 sky130_fd_sc_hd__nand2_1 _22210_ (.A(_11673_),
    .B(_12131_),
    .Y(_12133_));
 sky130_fd_sc_hd__a21oi_1 _22211_ (.A1(_11673_),
    .A2(_12131_),
    .B1(_11674_),
    .Y(_12134_));
 sky130_fd_sc_hd__o311a_1 _22212_ (.A1(_11178_),
    .A2(_11672_),
    .A3(_11676_),
    .B1(_12133_),
    .C1(_11675_),
    .X(_12135_));
 sky130_fd_sc_hd__o211ai_4 _22213_ (.A1(_11678_),
    .A2(_11672_),
    .B1(_11675_),
    .C1(_12133_),
    .Y(_12136_));
 sky130_fd_sc_hd__nand3_4 _22214_ (.A(_11673_),
    .B(_11675_),
    .C(_12131_),
    .Y(_12137_));
 sky130_fd_sc_hd__and4b_1 _22215_ (.A_N(_10227_),
    .B(_11673_),
    .C(_11675_),
    .D(_12131_),
    .X(_12138_));
 sky130_fd_sc_hd__nand4b_2 _22216_ (.A_N(_10227_),
    .B(_11673_),
    .C(_11675_),
    .D(_12131_),
    .Y(_12139_));
 sky130_fd_sc_hd__a2bb2oi_4 _22217_ (.A1_N(_10227_),
    .A2_N(_12137_),
    .B1(_11680_),
    .B2(_12134_),
    .Y(_12140_));
 sky130_fd_sc_hd__o21ai_1 _22218_ (.A1(_10227_),
    .A2(_12137_),
    .B1(_12136_),
    .Y(_12141_));
 sky130_fd_sc_hd__nand4_4 _22219_ (.A(_12125_),
    .B(_12128_),
    .C(_12136_),
    .D(_12139_),
    .Y(_12142_));
 sky130_fd_sc_hd__o21ai_4 _22220_ (.A1(_12124_),
    .A2(_12127_),
    .B1(_12141_),
    .Y(_12144_));
 sky130_fd_sc_hd__o221a_1 _22221_ (.A1(net302),
    .A2(_04019_),
    .B1(_12129_),
    .B2(_12140_),
    .C1(_12142_),
    .X(_12145_));
 sky130_fd_sc_hd__o221ai_4 _22222_ (.A1(net302),
    .A2(_04019_),
    .B1(_12129_),
    .B2(_12140_),
    .C1(_12142_),
    .Y(_12146_));
 sky130_fd_sc_hd__a31oi_4 _22223_ (.A1(_12144_),
    .A2(net277),
    .A3(_12142_),
    .B1(_12122_),
    .Y(_12147_));
 sky130_fd_sc_hd__o22a_4 _22224_ (.A1(_05228_),
    .A2(_05230_),
    .B1(_12122_),
    .B2(_12145_),
    .X(_12148_));
 sky130_fd_sc_hd__or3_2 _22225_ (.A(net296),
    .B(_05232_),
    .C(_12147_),
    .X(_12149_));
 sky130_fd_sc_hd__a31oi_1 _22226_ (.A1(_12144_),
    .A2(net277),
    .A3(_12142_),
    .B1(net232),
    .Y(_12150_));
 sky130_fd_sc_hd__o21ai_1 _22227_ (.A1(_06626_),
    .A2(_06627_),
    .B1(_12146_),
    .Y(_12151_));
 sky130_fd_sc_hd__a311oi_4 _22228_ (.A1(_12144_),
    .A2(net277),
    .A3(_12142_),
    .B1(net232),
    .C1(_12122_),
    .Y(_12152_));
 sky130_fd_sc_hd__nand3_2 _22229_ (.A(_12146_),
    .B(net234),
    .C(_12123_),
    .Y(_12153_));
 sky130_fd_sc_hd__a2bb2oi_2 _22230_ (.A1_N(_06622_),
    .A2_N(_06624_),
    .B1(_12123_),
    .B2(_12146_),
    .Y(_12155_));
 sky130_fd_sc_hd__o22ai_4 _22231_ (.A1(_06622_),
    .A2(_06624_),
    .B1(_12122_),
    .B2(_12145_),
    .Y(_12156_));
 sky130_fd_sc_hd__a21oi_1 _22232_ (.A1(_12123_),
    .A2(_12150_),
    .B1(_12155_),
    .Y(_12157_));
 sky130_fd_sc_hd__a31o_1 _22233_ (.A1(_11194_),
    .A2(_11685_),
    .A3(_11688_),
    .B1(_11689_),
    .X(_12158_));
 sky130_fd_sc_hd__a31oi_4 _22234_ (.A1(_11194_),
    .A2(_11685_),
    .A3(_11688_),
    .B1(_11689_),
    .Y(_12159_));
 sky130_fd_sc_hd__o21ai_4 _22235_ (.A1(_12152_),
    .A2(_12155_),
    .B1(_12159_),
    .Y(_12160_));
 sky130_fd_sc_hd__o211ai_4 _22236_ (.A1(_12122_),
    .A2(_12151_),
    .B1(_12158_),
    .C1(_12156_),
    .Y(_12161_));
 sky130_fd_sc_hd__o311a_1 _22237_ (.A1(_12152_),
    .A2(_12155_),
    .A3(_12159_),
    .B1(net272),
    .C1(_12160_),
    .X(_12162_));
 sky130_fd_sc_hd__nand3_2 _22238_ (.A(_12160_),
    .B(_12161_),
    .C(net272),
    .Y(_12163_));
 sky130_fd_sc_hd__a31oi_4 _22239_ (.A1(_12160_),
    .A2(_12161_),
    .A3(net272),
    .B1(_12148_),
    .Y(_12164_));
 sky130_fd_sc_hd__a31o_1 _22240_ (.A1(_12160_),
    .A2(_12161_),
    .A3(net272),
    .B1(_12148_),
    .X(_12166_));
 sky130_fd_sc_hd__a21oi_1 _22241_ (.A1(_11212_),
    .A2(_11228_),
    .B1(_11702_),
    .Y(_12167_));
 sky130_fd_sc_hd__a31oi_2 _22242_ (.A1(_11212_),
    .A2(_11228_),
    .A3(_11701_),
    .B1(_11702_),
    .Y(_12168_));
 sky130_fd_sc_hd__a31oi_2 _22243_ (.A1(_12160_),
    .A2(_12161_),
    .A3(net272),
    .B1(net251),
    .Y(_12169_));
 sky130_fd_sc_hd__a311oi_4 _22244_ (.A1(_12160_),
    .A2(_12161_),
    .A3(net272),
    .B1(net251),
    .C1(_12148_),
    .Y(_12170_));
 sky130_fd_sc_hd__o211ai_4 _22245_ (.A1(net272),
    .A2(_12147_),
    .B1(_06314_),
    .C1(_12163_),
    .Y(_12171_));
 sky130_fd_sc_hd__a2bb2oi_4 _22246_ (.A1_N(_06305_),
    .A2_N(_06307_),
    .B1(_12149_),
    .B2(_12163_),
    .Y(_12172_));
 sky130_fd_sc_hd__o22ai_2 _22247_ (.A1(net284),
    .A2(_06307_),
    .B1(_12148_),
    .B2(_12162_),
    .Y(_12173_));
 sky130_fd_sc_hd__a21oi_1 _22248_ (.A1(_12149_),
    .A2(_12169_),
    .B1(_12172_),
    .Y(_12174_));
 sky130_fd_sc_hd__nand3b_1 _22249_ (.A_N(_12168_),
    .B(_12171_),
    .C(_12173_),
    .Y(_12175_));
 sky130_fd_sc_hd__o22ai_1 _22250_ (.A1(_11700_),
    .A2(_12167_),
    .B1(_12170_),
    .B2(_12172_),
    .Y(_12177_));
 sky130_fd_sc_hd__nand3_1 _22251_ (.A(_12175_),
    .B(_12177_),
    .C(net245),
    .Y(_12178_));
 sky130_fd_sc_hd__or3_1 _22252_ (.A(net270),
    .B(_05483_),
    .C(_12164_),
    .X(_12179_));
 sky130_fd_sc_hd__o211ai_2 _22253_ (.A1(_11700_),
    .A2(_12167_),
    .B1(_12171_),
    .C1(_12173_),
    .Y(_12180_));
 sky130_fd_sc_hd__o21bai_2 _22254_ (.A1(_12170_),
    .A2(_12172_),
    .B1_N(_12168_),
    .Y(_12181_));
 sky130_fd_sc_hd__o211ai_2 _22255_ (.A1(net270),
    .A2(_05483_),
    .B1(_12180_),
    .C1(_12181_),
    .Y(_12182_));
 sky130_fd_sc_hd__o211ai_4 _22256_ (.A1(_12166_),
    .A2(net245),
    .B1(net253),
    .C1(_12178_),
    .Y(_12183_));
 sky130_fd_sc_hd__a31oi_2 _22257_ (.A1(_12180_),
    .A2(_12181_),
    .A3(net245),
    .B1(net253),
    .Y(_12184_));
 sky130_fd_sc_hd__o221a_1 _22258_ (.A1(_06011_),
    .A2(_06012_),
    .B1(_12164_),
    .B2(net245),
    .C1(_12182_),
    .X(_12185_));
 sky130_fd_sc_hd__o221ai_4 _22259_ (.A1(_06011_),
    .A2(_06012_),
    .B1(_12164_),
    .B2(net245),
    .C1(_12182_),
    .Y(_12186_));
 sky130_fd_sc_hd__a21oi_1 _22260_ (.A1(_11239_),
    .A2(_11723_),
    .B1(_11718_),
    .Y(_12188_));
 sky130_fd_sc_hd__a21o_1 _22261_ (.A1(_11239_),
    .A2(_11723_),
    .B1(_11718_),
    .X(_12189_));
 sky130_fd_sc_hd__a31oi_2 _22262_ (.A1(_11239_),
    .A2(_11722_),
    .A3(_11723_),
    .B1(_11718_),
    .Y(_12190_));
 sky130_fd_sc_hd__o2bb2ai_4 _22263_ (.A1_N(_12183_),
    .A2_N(_12186_),
    .B1(_12188_),
    .B2(_11721_),
    .Y(_12191_));
 sky130_fd_sc_hd__o2111ai_4 _22264_ (.A1(net261),
    .A2(_11716_),
    .B1(_12183_),
    .C1(_12186_),
    .D1(_12189_),
    .Y(_12192_));
 sky130_fd_sc_hd__nand3_4 _22265_ (.A(_12191_),
    .B(_12192_),
    .C(net242),
    .Y(_12193_));
 sky130_fd_sc_hd__o311a_2 _22266_ (.A1(net245),
    .A2(_12148_),
    .A3(_12162_),
    .B1(_12178_),
    .C1(_05754_),
    .X(_12194_));
 sky130_fd_sc_hd__inv_2 _22267_ (.A(_12194_),
    .Y(_12195_));
 sky130_fd_sc_hd__a31oi_4 _22268_ (.A1(_12191_),
    .A2(_12192_),
    .A3(net242),
    .B1(_12194_),
    .Y(_12196_));
 sky130_fd_sc_hd__a21oi_4 _22269_ (.A1(_12193_),
    .A2(_12195_),
    .B1(net240),
    .Y(_12197_));
 sky130_fd_sc_hd__or3_1 _22270_ (.A(_05990_),
    .B(_05992_),
    .C(_12196_),
    .X(_12199_));
 sky130_fd_sc_hd__a21oi_4 _22271_ (.A1(_12193_),
    .A2(_12195_),
    .B1(net263),
    .Y(_12200_));
 sky130_fd_sc_hd__a22o_2 _22272_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_12193_),
    .B2(_12195_),
    .X(_12201_));
 sky130_fd_sc_hd__and3_1 _22273_ (.A(_12193_),
    .B(_12195_),
    .C(net263),
    .X(_12202_));
 sky130_fd_sc_hd__a311o_4 _22274_ (.A1(_12191_),
    .A2(_12192_),
    .A3(net242),
    .B1(_12194_),
    .C1(net261),
    .X(_12203_));
 sky130_fd_sc_hd__and4_1 _22275_ (.A(_10291_),
    .B(_10294_),
    .C(_10765_),
    .D(_10767_),
    .X(_12204_));
 sky130_fd_sc_hd__o21a_1 _22276_ (.A1(net295),
    .A2(_11251_),
    .B1(_12204_),
    .X(_12205_));
 sky130_fd_sc_hd__o211a_1 _22277_ (.A1(_11235_),
    .A2(_11258_),
    .B1(_12204_),
    .C1(_11262_),
    .X(_12206_));
 sky130_fd_sc_hd__nand4_2 _22278_ (.A(_12204_),
    .B(_11740_),
    .C(_11262_),
    .D(_11260_),
    .Y(_12207_));
 sky130_fd_sc_hd__o2111ai_2 _22279_ (.A1(net294),
    .A2(_11252_),
    .B1(_11740_),
    .C1(_10307_),
    .D1(_12205_),
    .Y(_12208_));
 sky130_fd_sc_hd__o221ai_4 _22280_ (.A1(_11734_),
    .A2(net292),
    .B1(_12206_),
    .B2(_11750_),
    .C1(_12208_),
    .Y(_12210_));
 sky130_fd_sc_hd__o211a_1 _22281_ (.A1(_11746_),
    .A2(_11739_),
    .B1(_11741_),
    .C1(_12207_),
    .X(_12211_));
 sky130_fd_sc_hd__o211ai_4 _22282_ (.A1(_11746_),
    .A2(_11739_),
    .B1(_11741_),
    .C1(_12207_),
    .Y(_12212_));
 sky130_fd_sc_hd__nand4_1 _22283_ (.A(_12204_),
    .B(_11262_),
    .C(_11260_),
    .D(_10307_),
    .Y(_12213_));
 sky130_fd_sc_hd__o2111ai_4 _22284_ (.A1(net294),
    .A2(_11252_),
    .B1(_11740_),
    .C1(_11741_),
    .D1(_12205_),
    .Y(_12214_));
 sky130_fd_sc_hd__nand4_1 _22285_ (.A(_12206_),
    .B(_11741_),
    .C(_11740_),
    .D(_10307_),
    .Y(_12215_));
 sky130_fd_sc_hd__a41o_1 _22286_ (.A1(_10307_),
    .A2(_11740_),
    .A3(_11741_),
    .A4(_12206_),
    .B1(_12211_),
    .X(_12216_));
 sky130_fd_sc_hd__o221ai_4 _22287_ (.A1(_05507_),
    .A2(_11735_),
    .B1(_12200_),
    .B2(_12202_),
    .C1(_12210_),
    .Y(_12217_));
 sky130_fd_sc_hd__o2bb2ai_1 _22288_ (.A1_N(net263),
    .A2_N(_12196_),
    .B1(_12213_),
    .B2(_11742_),
    .Y(_12218_));
 sky130_fd_sc_hd__o211ai_4 _22289_ (.A1(_12214_),
    .A2(_10306_),
    .B1(_12203_),
    .C1(_12212_),
    .Y(_12219_));
 sky130_fd_sc_hd__o2111ai_4 _22290_ (.A1(_12214_),
    .A2(_10306_),
    .B1(_12203_),
    .C1(_12212_),
    .D1(_12201_),
    .Y(_12221_));
 sky130_fd_sc_hd__o311a_1 _22291_ (.A1(_12200_),
    .A2(_12218_),
    .A3(_12211_),
    .B1(net240),
    .C1(_12217_),
    .X(_12222_));
 sky130_fd_sc_hd__o221ai_4 _22292_ (.A1(_05990_),
    .A2(_05992_),
    .B1(_12200_),
    .B2(_12219_),
    .C1(_12217_),
    .Y(_12223_));
 sky130_fd_sc_hd__o22a_2 _22293_ (.A1(_06286_),
    .A2(_06288_),
    .B1(_12197_),
    .B2(_12222_),
    .X(_12224_));
 sky130_fd_sc_hd__a22o_1 _22294_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_12199_),
    .B2(_12223_),
    .X(_12225_));
 sky130_fd_sc_hd__a31o_1 _22295_ (.A1(net240),
    .A2(_12217_),
    .A3(_12221_),
    .B1(net292),
    .X(_12226_));
 sky130_fd_sc_hd__a311oi_4 _22296_ (.A1(net240),
    .A2(_12217_),
    .A3(_12221_),
    .B1(_12197_),
    .C1(net292),
    .Y(_12227_));
 sky130_fd_sc_hd__o211ai_2 _22297_ (.A1(net240),
    .A2(_12196_),
    .B1(net267),
    .C1(_12223_),
    .Y(_12228_));
 sky130_fd_sc_hd__a21oi_2 _22298_ (.A1(_12199_),
    .A2(_12223_),
    .B1(_05507_),
    .Y(_12229_));
 sky130_fd_sc_hd__o22ai_4 _22299_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_12197_),
    .B2(_12222_),
    .Y(_12230_));
 sky130_fd_sc_hd__o22a_1 _22300_ (.A1(_11736_),
    .A2(_11761_),
    .B1(_11764_),
    .B2(_11760_),
    .X(_12232_));
 sky130_fd_sc_hd__a21oi_2 _22301_ (.A1(_11760_),
    .A2(_11763_),
    .B1(_11764_),
    .Y(_12233_));
 sky130_fd_sc_hd__o21bai_4 _22302_ (.A1(_12227_),
    .A2(_12229_),
    .B1_N(_12232_),
    .Y(_12234_));
 sky130_fd_sc_hd__o211ai_4 _22303_ (.A1(_12197_),
    .A2(_12226_),
    .B1(_12232_),
    .C1(_12230_),
    .Y(_12235_));
 sky130_fd_sc_hd__o311a_1 _22304_ (.A1(_12227_),
    .A2(_12229_),
    .A3(_12233_),
    .B1(net213),
    .C1(_12234_),
    .X(_12236_));
 sky130_fd_sc_hd__nand3_1 _22305_ (.A(_12234_),
    .B(_12235_),
    .C(net213),
    .Y(_12237_));
 sky130_fd_sc_hd__a31oi_4 _22306_ (.A1(_12234_),
    .A2(_12235_),
    .A3(net213),
    .B1(_12224_),
    .Y(_12238_));
 sky130_fd_sc_hd__or4_2 _22307_ (.A(_06608_),
    .B(_06610_),
    .C(_12224_),
    .D(_12236_),
    .X(_12239_));
 sky130_fd_sc_hd__o221a_1 _22308_ (.A1(_02137_),
    .A2(_11286_),
    .B1(net299),
    .B2(_11776_),
    .C1(_11302_),
    .X(_12240_));
 sky130_fd_sc_hd__o211a_1 _22309_ (.A1(_02148_),
    .A2(_11285_),
    .B1(_11780_),
    .C1(_11784_),
    .X(_12241_));
 sky130_fd_sc_hd__a31oi_2 _22310_ (.A1(_11289_),
    .A2(_11302_),
    .A3(_11778_),
    .B1(_11779_),
    .Y(_12243_));
 sky130_fd_sc_hd__a311oi_4 _22311_ (.A1(_12234_),
    .A2(_12235_),
    .A3(net213),
    .B1(_12224_),
    .C1(net294),
    .Y(_12244_));
 sky130_fd_sc_hd__o211ai_2 _22312_ (.A1(_05246_),
    .A2(_05247_),
    .B1(_12225_),
    .C1(_12237_),
    .Y(_12245_));
 sky130_fd_sc_hd__a2bb2oi_2 _22313_ (.A1_N(net318),
    .A2_N(net316),
    .B1(_12225_),
    .B2(_12237_),
    .Y(_12246_));
 sky130_fd_sc_hd__o22ai_1 _22314_ (.A1(net318),
    .A2(net316),
    .B1(_12224_),
    .B2(_12236_),
    .Y(_12247_));
 sky130_fd_sc_hd__nor2_1 _22315_ (.A(_12244_),
    .B(_12246_),
    .Y(_12248_));
 sky130_fd_sc_hd__o211ai_1 _22316_ (.A1(_11779_),
    .A2(_12240_),
    .B1(_12245_),
    .C1(_12247_),
    .Y(_12249_));
 sky130_fd_sc_hd__o22ai_1 _22317_ (.A1(_11777_),
    .A2(_12241_),
    .B1(_12244_),
    .B2(_12246_),
    .Y(_12250_));
 sky130_fd_sc_hd__nand3_2 _22318_ (.A(_12249_),
    .B(_12250_),
    .C(net210),
    .Y(_12251_));
 sky130_fd_sc_hd__or3_1 _22319_ (.A(_06608_),
    .B(net237),
    .C(_12238_),
    .X(_12252_));
 sky130_fd_sc_hd__o21ai_1 _22320_ (.A1(net295),
    .A2(_12238_),
    .B1(_12243_),
    .Y(_12254_));
 sky130_fd_sc_hd__o22ai_2 _22321_ (.A1(_11779_),
    .A2(_12240_),
    .B1(_12244_),
    .B2(_12246_),
    .Y(_12255_));
 sky130_fd_sc_hd__o221ai_4 _22322_ (.A1(_06608_),
    .A2(_06610_),
    .B1(_12244_),
    .B2(_12254_),
    .C1(_12255_),
    .Y(_12256_));
 sky130_fd_sc_hd__o31a_4 _22323_ (.A1(_06608_),
    .A2(net237),
    .A3(_12238_),
    .B1(_12256_),
    .X(_12257_));
 sky130_fd_sc_hd__o311a_1 _22324_ (.A1(net210),
    .A2(_12224_),
    .A3(_12236_),
    .B1(_12251_),
    .C1(_04238_),
    .X(_12258_));
 sky130_fd_sc_hd__o211ai_4 _22325_ (.A1(net341),
    .A2(_04184_),
    .B1(_12239_),
    .C1(_12251_),
    .Y(_12259_));
 sky130_fd_sc_hd__and3_2 _22326_ (.A(_12256_),
    .B(net299),
    .C(_12252_),
    .X(_12260_));
 sky130_fd_sc_hd__nand3_2 _22327_ (.A(_12256_),
    .B(net299),
    .C(_12252_),
    .Y(_12261_));
 sky130_fd_sc_hd__a21oi_1 _22328_ (.A1(_02148_),
    .A2(_11790_),
    .B1(_11797_),
    .Y(_12262_));
 sky130_fd_sc_hd__o21bai_2 _22329_ (.A1(_11793_),
    .A2(_11798_),
    .B1_N(_11791_),
    .Y(_12263_));
 sky130_fd_sc_hd__a21oi_2 _22330_ (.A1(_12259_),
    .A2(_12261_),
    .B1(_12263_),
    .Y(_12265_));
 sky130_fd_sc_hd__o2bb2ai_1 _22331_ (.A1_N(_12259_),
    .A2_N(_12261_),
    .B1(_12262_),
    .B2(_11793_),
    .Y(_12266_));
 sky130_fd_sc_hd__o21ai_1 _22332_ (.A1(_11791_),
    .A2(_11806_),
    .B1(_12259_),
    .Y(_12267_));
 sky130_fd_sc_hd__a31o_2 _22333_ (.A1(_12259_),
    .A2(_12261_),
    .A3(_12263_),
    .B1(_06904_),
    .X(_12268_));
 sky130_fd_sc_hd__o221ai_4 _22334_ (.A1(_06899_),
    .A2(_06901_),
    .B1(_12260_),
    .B2(_12267_),
    .C1(_12266_),
    .Y(_12269_));
 sky130_fd_sc_hd__a211o_1 _22335_ (.A1(_12252_),
    .A2(_12256_),
    .B1(_06899_),
    .C1(_06901_),
    .X(_12270_));
 sky130_fd_sc_hd__o32a_2 _22336_ (.A1(net230),
    .A2(_06901_),
    .A3(_12257_),
    .B1(_12265_),
    .B2(_12268_),
    .X(_12271_));
 sky130_fd_sc_hd__o22ai_2 _22337_ (.A1(net208),
    .A2(_12257_),
    .B1(_12265_),
    .B2(_12268_),
    .Y(_12272_));
 sky130_fd_sc_hd__a21oi_4 _22338_ (.A1(_12269_),
    .A2(_12270_),
    .B1(_02137_),
    .Y(_12273_));
 sky130_fd_sc_hd__o21ai_2 _22339_ (.A1(_02049_),
    .A2(net343),
    .B1(_12272_),
    .Y(_12274_));
 sky130_fd_sc_hd__o221a_1 _22340_ (.A1(net208),
    .A2(_12257_),
    .B1(_12265_),
    .B2(_12268_),
    .C1(_02137_),
    .X(_12276_));
 sky130_fd_sc_hd__o221ai_4 _22341_ (.A1(net208),
    .A2(_12257_),
    .B1(_12265_),
    .B2(_12268_),
    .C1(_02137_),
    .Y(_12277_));
 sky130_fd_sc_hd__a22oi_2 _22342_ (.A1(_11957_),
    .A2(_11958_),
    .B1(_12274_),
    .B2(_12277_),
    .Y(_12278_));
 sky130_fd_sc_hd__o2bb2ai_2 _22343_ (.A1_N(_11957_),
    .A2_N(_11958_),
    .B1(_12273_),
    .B2(_12276_),
    .Y(_12279_));
 sky130_fd_sc_hd__nand3_1 _22344_ (.A(_11957_),
    .B(_11958_),
    .C(_12277_),
    .Y(_12280_));
 sky130_fd_sc_hd__nand4_4 _22345_ (.A(_11957_),
    .B(_11958_),
    .C(_12274_),
    .D(_12277_),
    .Y(_12281_));
 sky130_fd_sc_hd__o22ai_2 _22346_ (.A1(_07227_),
    .A2(_07229_),
    .B1(_12273_),
    .B2(_12280_),
    .Y(_12282_));
 sky130_fd_sc_hd__nand3_2 _22347_ (.A(net185),
    .B(_12279_),
    .C(_12281_),
    .Y(_12283_));
 sky130_fd_sc_hd__and3_2 _22348_ (.A(_07228_),
    .B(_07230_),
    .C(_12272_),
    .X(_12284_));
 sky130_fd_sc_hd__or3_2 _22349_ (.A(_07227_),
    .B(_07229_),
    .C(_12271_),
    .X(_12285_));
 sky130_fd_sc_hd__o22ai_4 _22350_ (.A1(net185),
    .A2(_12271_),
    .B1(_12278_),
    .B2(_12282_),
    .Y(_12287_));
 sky130_fd_sc_hd__and3_2 _22351_ (.A(_07545_),
    .B(_07547_),
    .C(_12287_),
    .X(_12288_));
 sky130_fd_sc_hd__a211o_1 _22352_ (.A1(_12283_),
    .A2(_12285_),
    .B1(_07544_),
    .C1(net184),
    .X(_12289_));
 sky130_fd_sc_hd__a31o_1 _22353_ (.A1(net185),
    .A2(_12279_),
    .A3(_12281_),
    .B1(_00251_),
    .X(_12290_));
 sky130_fd_sc_hd__a311oi_4 _22354_ (.A1(net185),
    .A2(_12279_),
    .A3(_12281_),
    .B1(_12284_),
    .C1(_00251_),
    .Y(_12291_));
 sky130_fd_sc_hd__nand3_2 _22355_ (.A(_12283_),
    .B(_12285_),
    .C(_00240_),
    .Y(_12292_));
 sky130_fd_sc_hd__a21oi_2 _22356_ (.A1(_12283_),
    .A2(_12285_),
    .B1(_00240_),
    .Y(_12293_));
 sky130_fd_sc_hd__o21ai_4 _22357_ (.A1(_00174_),
    .A2(net344),
    .B1(_12287_),
    .Y(_12294_));
 sky130_fd_sc_hd__a31o_1 _22358_ (.A1(_11348_),
    .A2(_11828_),
    .A3(_11833_),
    .B1(_11834_),
    .X(_12295_));
 sky130_fd_sc_hd__a21oi_4 _22359_ (.A1(_11831_),
    .A2(_11833_),
    .B1(_11834_),
    .Y(_12296_));
 sky130_fd_sc_hd__o21ai_4 _22360_ (.A1(_12291_),
    .A2(_12293_),
    .B1(_12296_),
    .Y(_12298_));
 sky130_fd_sc_hd__o211ai_4 _22361_ (.A1(_12284_),
    .A2(_12290_),
    .B1(_12295_),
    .C1(_12294_),
    .Y(_12299_));
 sky130_fd_sc_hd__o311a_1 _22362_ (.A1(_12291_),
    .A2(_12293_),
    .A3(_12296_),
    .B1(net163),
    .C1(_12298_),
    .X(_12300_));
 sky130_fd_sc_hd__nand3_2 _22363_ (.A(_12298_),
    .B(_12299_),
    .C(net163),
    .Y(_12301_));
 sky130_fd_sc_hd__a31oi_4 _22364_ (.A1(_12298_),
    .A2(_12299_),
    .A3(net163),
    .B1(_12288_),
    .Y(_12302_));
 sky130_fd_sc_hd__a31o_1 _22365_ (.A1(_12298_),
    .A2(_12299_),
    .A3(net163),
    .B1(_12288_),
    .X(_12303_));
 sky130_fd_sc_hd__o311a_1 _22366_ (.A1(net365),
    .A2(net362),
    .A3(_11358_),
    .B1(_11371_),
    .C1(_11848_),
    .X(_12304_));
 sky130_fd_sc_hd__o211a_1 _22367_ (.A1(_11363_),
    .A2(_11365_),
    .B1(_11368_),
    .C1(_11849_),
    .X(_12305_));
 sky130_fd_sc_hd__a21o_1 _22368_ (.A1(_11849_),
    .A2(_11852_),
    .B1(_11846_),
    .X(_12306_));
 sky130_fd_sc_hd__a311oi_4 _22369_ (.A1(_12298_),
    .A2(_12299_),
    .A3(net163),
    .B1(_12288_),
    .C1(_12899_),
    .Y(_12307_));
 sky130_fd_sc_hd__o211ai_4 _22370_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_12289_),
    .C1(_12301_),
    .Y(_12309_));
 sky130_fd_sc_hd__a2bb2oi_2 _22371_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_12289_),
    .B2(_12301_),
    .Y(_12310_));
 sky130_fd_sc_hd__a2bb2o_1 _22372_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_12289_),
    .B2(_12301_),
    .X(_12311_));
 sky130_fd_sc_hd__o211ai_1 _22373_ (.A1(_11850_),
    .A2(_12304_),
    .B1(_12309_),
    .C1(_12311_),
    .Y(_12312_));
 sky130_fd_sc_hd__o22ai_1 _22374_ (.A1(_11846_),
    .A2(_12305_),
    .B1(_12307_),
    .B2(_12310_),
    .Y(_12313_));
 sky130_fd_sc_hd__nand3_2 _22375_ (.A(_12312_),
    .B(_12313_),
    .C(net160),
    .Y(_12314_));
 sky130_fd_sc_hd__and3_1 _22376_ (.A(_07913_),
    .B(_07915_),
    .C(_12303_),
    .X(_12315_));
 sky130_fd_sc_hd__or3_1 _22377_ (.A(_07912_),
    .B(_07914_),
    .C(_12302_),
    .X(_12316_));
 sky130_fd_sc_hd__o21ai_1 _22378_ (.A1(_12888_),
    .A2(_12302_),
    .B1(_12306_),
    .Y(_12317_));
 sky130_fd_sc_hd__o211ai_2 _22379_ (.A1(_11846_),
    .A2(_12305_),
    .B1(_12309_),
    .C1(_12311_),
    .Y(_12318_));
 sky130_fd_sc_hd__o22ai_4 _22380_ (.A1(_11850_),
    .A2(_12304_),
    .B1(_12307_),
    .B2(_12310_),
    .Y(_12320_));
 sky130_fd_sc_hd__o221ai_4 _22381_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_12307_),
    .B2(_12317_),
    .C1(_12320_),
    .Y(_12321_));
 sky130_fd_sc_hd__a31oi_4 _22382_ (.A1(_12318_),
    .A2(_12320_),
    .A3(net160),
    .B1(_12315_),
    .Y(_12322_));
 sky130_fd_sc_hd__a2bb2oi_1 _22383_ (.A1_N(_11210_),
    .A2_N(_11232_),
    .B1(_12316_),
    .B2(_12321_),
    .Y(_12323_));
 sky130_fd_sc_hd__o211ai_4 _22384_ (.A1(_12303_),
    .A2(net160),
    .B1(_11309_),
    .C1(_12314_),
    .Y(_12324_));
 sky130_fd_sc_hd__and3_1 _22385_ (.A(_12321_),
    .B(_11298_),
    .C(_12316_),
    .X(_12325_));
 sky130_fd_sc_hd__o211ai_4 _22386_ (.A1(net160),
    .A2(_12302_),
    .B1(_11298_),
    .C1(_12321_),
    .Y(_12326_));
 sky130_fd_sc_hd__o311a_1 _22387_ (.A1(_10881_),
    .A2(_11379_),
    .A3(_11381_),
    .B1(_11384_),
    .C1(_11860_),
    .X(_12327_));
 sky130_fd_sc_hd__o21ai_2 _22388_ (.A1(_11861_),
    .A2(_11864_),
    .B1(_11860_),
    .Y(_12328_));
 sky130_fd_sc_hd__a21oi_4 _22389_ (.A1(_12324_),
    .A2(_12326_),
    .B1(_12328_),
    .Y(_12329_));
 sky130_fd_sc_hd__o2bb2ai_1 _22390_ (.A1_N(_12324_),
    .A2_N(_12326_),
    .B1(_12327_),
    .B2(_11861_),
    .Y(_12331_));
 sky130_fd_sc_hd__nand3_1 _22391_ (.A(_12324_),
    .B(_12326_),
    .C(_12328_),
    .Y(_12332_));
 sky130_fd_sc_hd__a31o_2 _22392_ (.A1(_12324_),
    .A2(_12326_),
    .A3(_12328_),
    .B1(_08301_),
    .X(_12333_));
 sky130_fd_sc_hd__nand3_1 _22393_ (.A(_12331_),
    .B(_12332_),
    .C(_08300_),
    .Y(_12334_));
 sky130_fd_sc_hd__o311a_1 _22394_ (.A1(net160),
    .A2(_12288_),
    .A3(_12300_),
    .B1(_12314_),
    .C1(_08301_),
    .X(_12335_));
 sky130_fd_sc_hd__or3_1 _22395_ (.A(net180),
    .B(_08298_),
    .C(_12322_),
    .X(_12336_));
 sky130_fd_sc_hd__o32a_2 _22396_ (.A1(net180),
    .A2(_08298_),
    .A3(_12322_),
    .B1(_12329_),
    .B2(_12333_),
    .X(_12337_));
 sky130_fd_sc_hd__o22ai_2 _22397_ (.A1(_08300_),
    .A2(_12322_),
    .B1(_12329_),
    .B2(_12333_),
    .Y(_12338_));
 sky130_fd_sc_hd__a22oi_4 _22398_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_12334_),
    .B2(_12336_),
    .Y(_12339_));
 sky130_fd_sc_hd__o21ai_2 _22399_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_12338_),
    .Y(_12340_));
 sky130_fd_sc_hd__o22ai_1 _22400_ (.A1(net365),
    .A2(net362),
    .B1(_12329_),
    .B2(_12333_),
    .Y(_12342_));
 sky130_fd_sc_hd__o221a_1 _22401_ (.A1(_08300_),
    .A2(_12322_),
    .B1(_12329_),
    .B2(_12333_),
    .C1(_10015_),
    .X(_12343_));
 sky130_fd_sc_hd__o221ai_4 _22402_ (.A1(_08300_),
    .A2(_12322_),
    .B1(_12329_),
    .B2(_12333_),
    .C1(_10015_),
    .Y(_12344_));
 sky130_fd_sc_hd__a21oi_4 _22403_ (.A1(_12340_),
    .A2(_12344_),
    .B1(_11951_),
    .Y(_12345_));
 sky130_fd_sc_hd__o21bai_1 _22404_ (.A1(_12339_),
    .A2(_12343_),
    .B1_N(_11951_),
    .Y(_12346_));
 sky130_fd_sc_hd__o2bb2ai_2 _22405_ (.A1_N(_11882_),
    .A2_N(_11950_),
    .B1(_12335_),
    .B2(_12342_),
    .Y(_12347_));
 sky130_fd_sc_hd__o22ai_4 _22406_ (.A1(net158),
    .A2(_08712_),
    .B1(_12339_),
    .B2(_12347_),
    .Y(_12348_));
 sky130_fd_sc_hd__o211ai_2 _22407_ (.A1(_12339_),
    .A2(_12347_),
    .B1(_08714_),
    .C1(_12346_),
    .Y(_12349_));
 sky130_fd_sc_hd__or3_2 _22408_ (.A(net158),
    .B(_08712_),
    .C(_12337_),
    .X(_12350_));
 sky130_fd_sc_hd__o21ai_4 _22409_ (.A1(_12345_),
    .A2(_12348_),
    .B1(_12350_),
    .Y(_12351_));
 sky130_fd_sc_hd__a32oi_4 _22410_ (.A1(_11890_),
    .A2(_07877_),
    .A3(_07855_),
    .B1(_11896_),
    .B2(_11893_),
    .Y(_12353_));
 sky130_fd_sc_hd__a32o_1 _22411_ (.A1(_11890_),
    .A2(_07877_),
    .A3(_07855_),
    .B1(_11896_),
    .B2(_11893_),
    .X(_12354_));
 sky130_fd_sc_hd__o221a_1 _22412_ (.A1(_08714_),
    .A2(_12337_),
    .B1(_12345_),
    .B2(_12348_),
    .C1(_08907_),
    .X(_12355_));
 sky130_fd_sc_hd__o221ai_4 _22413_ (.A1(_08714_),
    .A2(_12337_),
    .B1(_12345_),
    .B2(_12348_),
    .C1(_08907_),
    .Y(_12356_));
 sky130_fd_sc_hd__a21oi_1 _22414_ (.A1(_12349_),
    .A2(_12350_),
    .B1(_08907_),
    .Y(_12357_));
 sky130_fd_sc_hd__o21ai_2 _22415_ (.A1(_08819_),
    .A2(_08841_),
    .B1(_12351_),
    .Y(_12358_));
 sky130_fd_sc_hd__nand3_1 _22416_ (.A(_12354_),
    .B(_12356_),
    .C(_12358_),
    .Y(_12359_));
 sky130_fd_sc_hd__o21ai_1 _22417_ (.A1(_12355_),
    .A2(_12357_),
    .B1(_12353_),
    .Y(_12360_));
 sky130_fd_sc_hd__nand3_1 _22418_ (.A(_12358_),
    .B(_12353_),
    .C(_12356_),
    .Y(_12361_));
 sky130_fd_sc_hd__o21ai_1 _22419_ (.A1(_12355_),
    .A2(_12357_),
    .B1(_12354_),
    .Y(_12362_));
 sky130_fd_sc_hd__o211ai_4 _22420_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_12361_),
    .C1(_12362_),
    .Y(_12364_));
 sky130_fd_sc_hd__a211o_1 _22421_ (.A1(_12349_),
    .A2(_12350_),
    .B1(_09120_),
    .C1(_09121_),
    .X(_12365_));
 sky130_fd_sc_hd__o211ai_2 _22422_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_12359_),
    .C1(_12360_),
    .Y(_12366_));
 sky130_fd_sc_hd__o31a_2 _22423_ (.A1(_09120_),
    .A2(_09121_),
    .A3(_12351_),
    .B1(_12364_),
    .X(_12367_));
 sky130_fd_sc_hd__o211a_2 _22424_ (.A1(_09125_),
    .A2(_12351_),
    .B1(_12364_),
    .C1(_07899_),
    .X(_12368_));
 sky130_fd_sc_hd__o211ai_4 _22425_ (.A1(_09125_),
    .A2(_12351_),
    .B1(_12364_),
    .C1(_07899_),
    .Y(_12369_));
 sky130_fd_sc_hd__o211ai_4 _22426_ (.A1(net368),
    .A2(_07866_),
    .B1(_12365_),
    .C1(_12366_),
    .Y(_12370_));
 sky130_fd_sc_hd__o221a_1 _22427_ (.A1(_11422_),
    .A2(_06332_),
    .B1(_07033_),
    .B2(_11901_),
    .C1(_11431_),
    .X(_12371_));
 sky130_fd_sc_hd__o22a_1 _22428_ (.A1(_11900_),
    .A2(_11905_),
    .B1(_11424_),
    .B2(_11429_),
    .X(_12372_));
 sky130_fd_sc_hd__o21ai_1 _22429_ (.A1(_11904_),
    .A2(_11906_),
    .B1(_11908_),
    .Y(_12373_));
 sky130_fd_sc_hd__o2111ai_4 _22430_ (.A1(_11904_),
    .A2(_11906_),
    .B1(_11908_),
    .C1(_12369_),
    .D1(_12370_),
    .Y(_12375_));
 sky130_fd_sc_hd__o2bb2ai_1 _22431_ (.A1_N(_12369_),
    .A2_N(_12370_),
    .B1(_12372_),
    .B2(_11907_),
    .Y(_12376_));
 sky130_fd_sc_hd__o2111ai_4 _22432_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .C1(_12375_),
    .D1(_12376_),
    .Y(_12377_));
 sky130_fd_sc_hd__a211o_1 _22433_ (.A1(_12365_),
    .A2(_12366_),
    .B1(_09553_),
    .C1(net155),
    .X(_12378_));
 sky130_fd_sc_hd__o2bb2ai_1 _22434_ (.A1_N(_12369_),
    .A2_N(_12370_),
    .B1(_12371_),
    .B2(_11906_),
    .Y(_12379_));
 sky130_fd_sc_hd__o22a_1 _22435_ (.A1(_11907_),
    .A2(_12372_),
    .B1(_07899_),
    .B2(_12367_),
    .X(_12380_));
 sky130_fd_sc_hd__o21ai_2 _22436_ (.A1(_11907_),
    .A2(_12372_),
    .B1(_12370_),
    .Y(_12381_));
 sky130_fd_sc_hd__o211ai_2 _22437_ (.A1(_12381_),
    .A2(_12368_),
    .B1(net143),
    .C1(_12379_),
    .Y(_12382_));
 sky130_fd_sc_hd__nand2_1 _22438_ (.A(_12378_),
    .B(_12382_),
    .Y(_12383_));
 sky130_fd_sc_hd__a21oi_2 _22439_ (.A1(_11916_),
    .A2(_11917_),
    .B1(_11914_),
    .Y(_12384_));
 sky130_fd_sc_hd__a21o_1 _22440_ (.A1(_11916_),
    .A2(_11917_),
    .B1(_11914_),
    .X(_12386_));
 sky130_fd_sc_hd__and3_1 _22441_ (.A(_12382_),
    .B(_07033_),
    .C(_12378_),
    .X(_12387_));
 sky130_fd_sc_hd__o211ai_2 _22442_ (.A1(_06989_),
    .A2(net375),
    .B1(_12378_),
    .C1(_12382_),
    .Y(_12388_));
 sky130_fd_sc_hd__o211a_1 _22443_ (.A1(_12367_),
    .A2(net143),
    .B1(_07044_),
    .C1(_12377_),
    .X(_12389_));
 sky130_fd_sc_hd__o2111ai_4 _22444_ (.A1(_12367_),
    .A2(net143),
    .B1(_07022_),
    .C1(net376),
    .D1(_12377_),
    .Y(_12390_));
 sky130_fd_sc_hd__a21oi_1 _22445_ (.A1(_12388_),
    .A2(_12390_),
    .B1(_12384_),
    .Y(_12391_));
 sky130_fd_sc_hd__a31o_1 _22446_ (.A1(_12388_),
    .A2(_12390_),
    .A3(_12384_),
    .B1(_09578_),
    .X(_12392_));
 sky130_fd_sc_hd__o22a_2 _22447_ (.A1(_09579_),
    .A2(_12383_),
    .B1(_12391_),
    .B2(_12392_),
    .X(_12393_));
 sky130_fd_sc_hd__o221a_1 _22448_ (.A1(_09579_),
    .A2(_12383_),
    .B1(_12391_),
    .B2(_12392_),
    .C1(_06343_),
    .X(_12394_));
 sky130_fd_sc_hd__o21ai_2 _22449_ (.A1(net394),
    .A2(_06267_),
    .B1(_12393_),
    .Y(_12395_));
 sky130_fd_sc_hd__a21oi_1 _22450_ (.A1(_06300_),
    .A2(_06321_),
    .B1(_12393_),
    .Y(_12397_));
 sky130_fd_sc_hd__o21ba_1 _22451_ (.A1(_11926_),
    .A2(_11922_),
    .B1_N(_11925_),
    .X(_12398_));
 sky130_fd_sc_hd__o21bai_1 _22452_ (.A1(_12394_),
    .A2(_12397_),
    .B1_N(_12398_),
    .Y(_12399_));
 sky130_fd_sc_hd__o21ai_4 _22453_ (.A1(_06343_),
    .A2(_12393_),
    .B1(_12398_),
    .Y(_12400_));
 sky130_fd_sc_hd__o221ai_4 _22454_ (.A1(_10474_),
    .A2(net138),
    .B1(_12394_),
    .B2(_12400_),
    .C1(_12399_),
    .Y(_12401_));
 sky130_fd_sc_hd__o21ai_1 _22455_ (.A1(_10477_),
    .A2(_10478_),
    .B1(_12393_),
    .Y(_12402_));
 sky130_fd_sc_hd__o21ai_2 _22456_ (.A1(_11931_),
    .A2(_11929_),
    .B1(_11930_),
    .Y(_12403_));
 sky130_fd_sc_hd__o21ai_2 _22457_ (.A1(_05807_),
    .A2(_05829_),
    .B1(_12403_),
    .Y(_12404_));
 sky130_fd_sc_hd__o311ai_2 _22458_ (.A1(_05807_),
    .A2(_05829_),
    .A3(_12403_),
    .B1(_12404_),
    .C1(_10954_),
    .Y(_12405_));
 sky130_fd_sc_hd__a21oi_1 _22459_ (.A1(_12401_),
    .A2(_12402_),
    .B1(_12405_),
    .Y(_12406_));
 sky130_fd_sc_hd__a31oi_1 _22460_ (.A1(_12401_),
    .A2(_12402_),
    .A3(_12405_),
    .B1(_12406_),
    .Y(_12408_));
 sky130_fd_sc_hd__o21ai_1 _22461_ (.A1(_05250_),
    .A2(_11936_),
    .B1(_11940_),
    .Y(_12409_));
 sky130_fd_sc_hd__o21ai_1 _22462_ (.A1(_05447_),
    .A2(_05469_),
    .B1(_12409_),
    .Y(_12410_));
 sky130_fd_sc_hd__a21o_1 _22463_ (.A1(_05512_),
    .A2(net396),
    .B1(_12409_),
    .X(_12411_));
 sky130_fd_sc_hd__and4_1 _22464_ (.A(_11465_),
    .B(_12411_),
    .C(_12408_),
    .D(_12410_),
    .X(_12412_));
 sky130_fd_sc_hd__a31oi_1 _22465_ (.A1(_11465_),
    .A2(_12410_),
    .A3(_12411_),
    .B1(_12408_),
    .Y(_12413_));
 sky130_fd_sc_hd__or2_1 _22466_ (.A(_12412_),
    .B(_12413_),
    .X(_12414_));
 sky130_fd_sc_hd__o22a_1 _22467_ (.A1(net407),
    .A2(_05218_),
    .B1(_03289_),
    .B2(_11942_),
    .X(_12415_));
 sky130_fd_sc_hd__o21a_1 _22468_ (.A1(_11944_),
    .A2(_12415_),
    .B1(_12414_),
    .X(_12416_));
 sky130_fd_sc_hd__xnor2_1 _22469_ (.A(_11949_),
    .B(_12416_),
    .Y(net90));
 sky130_fd_sc_hd__nor3b_2 _22470_ (.A(_11468_),
    .B(_11945_),
    .C_N(_12416_),
    .Y(_12418_));
 sky130_fd_sc_hd__o31a_2 _22471_ (.A1(_11470_),
    .A2(_11961_),
    .A3(_11965_),
    .B1(_05403_),
    .X(_12419_));
 sky130_fd_sc_hd__o311a_1 _22472_ (.A1(_11470_),
    .A2(_11961_),
    .A3(_11965_),
    .B1(_05731_),
    .C1(_05403_),
    .X(_12420_));
 sky130_fd_sc_hd__or3b_1 _22473_ (.A(_10965_),
    .B(_10967_),
    .C_N(_12419_),
    .X(_12421_));
 sky130_fd_sc_hd__xor2_2 _22474_ (.A(_10970_),
    .B(_12419_),
    .X(_12422_));
 sky130_fd_sc_hd__o21bai_2 _22475_ (.A1(_11972_),
    .A2(_11979_),
    .B1_N(_12422_),
    .Y(_12423_));
 sky130_fd_sc_hd__o211ai_4 _22476_ (.A1(_11976_),
    .A2(_11977_),
    .B1(_12422_),
    .C1(_11973_),
    .Y(_12424_));
 sky130_fd_sc_hd__nor2_2 _22477_ (.A(net358),
    .B(_12419_),
    .Y(_12425_));
 sky130_fd_sc_hd__a21oi_4 _22478_ (.A1(_12423_),
    .A2(_12424_),
    .B1(_05731_),
    .Y(_12426_));
 sky130_fd_sc_hd__a31oi_2 _22479_ (.A1(_12423_),
    .A2(_12424_),
    .A3(net358),
    .B1(_12420_),
    .Y(_12427_));
 sky130_fd_sc_hd__or4_2 _22480_ (.A(_06793_),
    .B(_06815_),
    .C(_12425_),
    .D(_12426_),
    .X(_12429_));
 sky130_fd_sc_hd__or4_2 _22481_ (.A(_10489_),
    .B(_10490_),
    .C(_12425_),
    .D(_12426_),
    .X(_12430_));
 sky130_fd_sc_hd__o21ai_2 _22482_ (.A1(_10489_),
    .A2(_10490_),
    .B1(_12427_),
    .Y(_12431_));
 sky130_fd_sc_hd__o41a_1 _22483_ (.A1(_10489_),
    .A2(_10490_),
    .A3(_12425_),
    .A4(_12426_),
    .B1(_12431_),
    .X(_12432_));
 sky130_fd_sc_hd__o41ai_4 _22484_ (.A1(_10489_),
    .A2(_10490_),
    .A3(_12425_),
    .A4(_12426_),
    .B1(_12431_),
    .Y(_12433_));
 sky130_fd_sc_hd__a22oi_4 _22485_ (.A1(net151),
    .A2(_11983_),
    .B1(_11991_),
    .B2(_12001_),
    .Y(_12434_));
 sky130_fd_sc_hd__o221ai_4 _22486_ (.A1(_10026_),
    .A2(_11982_),
    .B1(_11992_),
    .B2(_12002_),
    .C1(_12433_),
    .Y(_12435_));
 sky130_fd_sc_hd__o21ai_4 _22487_ (.A1(_11986_),
    .A2(_12004_),
    .B1(_12432_),
    .Y(_12436_));
 sky130_fd_sc_hd__o211ai_4 _22488_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_12435_),
    .C1(_12436_),
    .Y(_12437_));
 sky130_fd_sc_hd__o31a_4 _22489_ (.A1(net357),
    .A2(_12425_),
    .A3(_12426_),
    .B1(_12437_),
    .X(_12438_));
 sky130_fd_sc_hd__a2bb2oi_1 _22490_ (.A1_N(_10021_),
    .A2_N(_10022_),
    .B1(_12429_),
    .B2(_12437_),
    .Y(_12440_));
 sky130_fd_sc_hd__a2bb2o_1 _22491_ (.A1_N(_10021_),
    .A2_N(_10022_),
    .B1(_12429_),
    .B2(_12437_),
    .X(_12441_));
 sky130_fd_sc_hd__a31oi_2 _22492_ (.A1(_12436_),
    .A2(net357),
    .A3(_12435_),
    .B1(net151),
    .Y(_12442_));
 sky130_fd_sc_hd__and3_1 _22493_ (.A(_12437_),
    .B(_10026_),
    .C(_12429_),
    .X(_12443_));
 sky130_fd_sc_hd__o21ai_1 _22494_ (.A1(net357),
    .A2(_12427_),
    .B1(_12442_),
    .Y(_12444_));
 sky130_fd_sc_hd__a21oi_2 _22495_ (.A1(_12429_),
    .A2(_12442_),
    .B1(_12440_),
    .Y(_12445_));
 sky130_fd_sc_hd__nand2_4 _22496_ (.A(_12441_),
    .B(_12444_),
    .Y(_12446_));
 sky130_fd_sc_hd__and3_1 _22497_ (.A(_11043_),
    .B(_11045_),
    .C(_10566_),
    .X(_12447_));
 sky130_fd_sc_hd__nand3_1 _22498_ (.A(_11043_),
    .B(_11045_),
    .C(_10566_),
    .Y(_12448_));
 sky130_fd_sc_hd__nor3_1 _22499_ (.A(_11533_),
    .B(_11534_),
    .C(_12448_),
    .Y(_12449_));
 sky130_fd_sc_hd__a21oi_2 _22500_ (.A1(_12449_),
    .A2(_12014_),
    .B1(_12015_),
    .Y(_12451_));
 sky130_fd_sc_hd__nand2_1 _22501_ (.A(_12017_),
    .B(_12451_),
    .Y(_12452_));
 sky130_fd_sc_hd__nand4_4 _22502_ (.A(_12014_),
    .B(_12447_),
    .C(_10573_),
    .D(_11536_),
    .Y(_12453_));
 sky130_fd_sc_hd__a21o_1 _22503_ (.A1(_09595_),
    .A2(_12008_),
    .B1(_12453_),
    .X(_12454_));
 sky130_fd_sc_hd__a2bb2oi_1 _22504_ (.A1_N(_12453_),
    .A2_N(_12015_),
    .B1(_12451_),
    .B2(_12017_),
    .Y(_12455_));
 sky130_fd_sc_hd__o2bb2ai_4 _22505_ (.A1_N(_12451_),
    .A2_N(_12017_),
    .B1(_12015_),
    .B2(_12453_),
    .Y(_12456_));
 sky130_fd_sc_hd__a21oi_2 _22506_ (.A1(_12452_),
    .A2(_12454_),
    .B1(_12445_),
    .Y(_12457_));
 sky130_fd_sc_hd__o21ai_2 _22507_ (.A1(_12440_),
    .A2(_12443_),
    .B1(_12456_),
    .Y(_12458_));
 sky130_fd_sc_hd__o211ai_2 _22508_ (.A1(_12015_),
    .A2(_12453_),
    .B1(_12452_),
    .C1(_12445_),
    .Y(_12459_));
 sky130_fd_sc_hd__o22ai_4 _22509_ (.A1(net374),
    .A2(_07702_),
    .B1(_12446_),
    .B2(_12456_),
    .Y(_12460_));
 sky130_fd_sc_hd__o221ai_4 _22510_ (.A1(net374),
    .A2(_07702_),
    .B1(_12446_),
    .B2(_12456_),
    .C1(_12458_),
    .Y(_12462_));
 sky130_fd_sc_hd__a21oi_1 _22511_ (.A1(_12429_),
    .A2(_12437_),
    .B1(net354),
    .Y(_12463_));
 sky130_fd_sc_hd__or3_1 _22512_ (.A(net374),
    .B(_07702_),
    .C(_12438_),
    .X(_12464_));
 sky130_fd_sc_hd__o22ai_4 _22513_ (.A1(net354),
    .A2(_12438_),
    .B1(_12457_),
    .B2(_12460_),
    .Y(_12465_));
 sky130_fd_sc_hd__and3_2 _22514_ (.A(_08689_),
    .B(_08711_),
    .C(_12465_),
    .X(_12466_));
 sky130_fd_sc_hd__inv_2 _22515_ (.A(_12466_),
    .Y(_12467_));
 sky130_fd_sc_hd__a221oi_2 _22516_ (.A1(net173),
    .A2(_12021_),
    .B1(_11553_),
    .B2(_11549_),
    .C1(_11546_),
    .Y(_12468_));
 sky130_fd_sc_hd__o221ai_1 _22517_ (.A1(net174),
    .A2(_12020_),
    .B1(_11548_),
    .B2(_11554_),
    .C1(_11547_),
    .Y(_12469_));
 sky130_fd_sc_hd__a31oi_2 _22518_ (.A1(_11547_),
    .A2(_11555_),
    .A3(_12024_),
    .B1(_12026_),
    .Y(_12470_));
 sky130_fd_sc_hd__o21ai_1 _22519_ (.A1(net173),
    .A2(_12021_),
    .B1(_12469_),
    .Y(_12471_));
 sky130_fd_sc_hd__a311oi_4 _22520_ (.A1(_12458_),
    .A2(_12459_),
    .A3(net354),
    .B1(_12463_),
    .C1(_09595_),
    .Y(_12473_));
 sky130_fd_sc_hd__o221ai_4 _22521_ (.A1(net354),
    .A2(_12438_),
    .B1(_12457_),
    .B2(_12460_),
    .C1(net172),
    .Y(_12474_));
 sky130_fd_sc_hd__a22oi_4 _22522_ (.A1(_09589_),
    .A2(_09591_),
    .B1(_12462_),
    .B2(_12464_),
    .Y(_12475_));
 sky130_fd_sc_hd__o21ai_4 _22523_ (.A1(_09588_),
    .A2(net187),
    .B1(_12465_),
    .Y(_12476_));
 sky130_fd_sc_hd__nand3_4 _22524_ (.A(_12470_),
    .B(_12474_),
    .C(_12476_),
    .Y(_12477_));
 sky130_fd_sc_hd__o22ai_4 _22525_ (.A1(_12026_),
    .A2(_12468_),
    .B1(_12473_),
    .B2(_12475_),
    .Y(_12478_));
 sky130_fd_sc_hd__o211ai_2 _22526_ (.A1(_08678_),
    .A2(_08700_),
    .B1(_12477_),
    .C1(_12478_),
    .Y(_12479_));
 sky130_fd_sc_hd__a31oi_4 _22527_ (.A1(_12477_),
    .A2(_12478_),
    .A3(net338),
    .B1(_12466_),
    .Y(_12480_));
 sky130_fd_sc_hd__a31o_1 _22528_ (.A1(_12477_),
    .A2(_12478_),
    .A3(net338),
    .B1(_12466_),
    .X(_12481_));
 sky130_fd_sc_hd__o31ai_2 _22529_ (.A1(_11566_),
    .A2(_12043_),
    .A3(_12046_),
    .B1(_12042_),
    .Y(_12482_));
 sky130_fd_sc_hd__a311oi_4 _22530_ (.A1(_12477_),
    .A2(_12478_),
    .A3(net338),
    .B1(net173),
    .C1(_12466_),
    .Y(_12484_));
 sky130_fd_sc_hd__a311o_2 _22531_ (.A1(_12477_),
    .A2(_12478_),
    .A3(net338),
    .B1(net173),
    .C1(_12466_),
    .X(_12485_));
 sky130_fd_sc_hd__a2bb2oi_4 _22532_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_12467_),
    .B2(_12479_),
    .Y(_12486_));
 sky130_fd_sc_hd__a2bb2o_1 _22533_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_12467_),
    .B2(_12479_),
    .X(_12487_));
 sky130_fd_sc_hd__nand3_2 _22534_ (.A(_12482_),
    .B(_12485_),
    .C(_12487_),
    .Y(_12488_));
 sky130_fd_sc_hd__o221ai_4 _22535_ (.A1(net177),
    .A2(_12039_),
    .B1(_12484_),
    .B2(_12486_),
    .C1(_12049_),
    .Y(_12489_));
 sky130_fd_sc_hd__and3_1 _22536_ (.A(_09796_),
    .B(_09818_),
    .C(_12481_),
    .X(_12490_));
 sky130_fd_sc_hd__or3_2 _22537_ (.A(net351),
    .B(_09807_),
    .C(_12480_),
    .X(_12491_));
 sky130_fd_sc_hd__nand3_2 _22538_ (.A(_12488_),
    .B(_12489_),
    .C(net335),
    .Y(_12492_));
 sky130_fd_sc_hd__a31o_1 _22539_ (.A1(_12488_),
    .A2(_12489_),
    .A3(net335),
    .B1(_12490_),
    .X(_12493_));
 sky130_fd_sc_hd__a31oi_2 _22540_ (.A1(_12488_),
    .A2(_12489_),
    .A3(net335),
    .B1(_12490_),
    .Y(_12495_));
 sky130_fd_sc_hd__o311a_1 _22541_ (.A1(net351),
    .A2(_09807_),
    .A3(_12480_),
    .B1(_12492_),
    .C1(_11079_),
    .X(_12496_));
 sky130_fd_sc_hd__a21oi_2 _22542_ (.A1(_12491_),
    .A2(_12492_),
    .B1(net177),
    .Y(_12497_));
 sky130_fd_sc_hd__a22o_2 _22543_ (.A1(_08725_),
    .A2(_08727_),
    .B1(_12491_),
    .B2(_12492_),
    .X(_12498_));
 sky130_fd_sc_hd__o211a_2 _22544_ (.A1(net335),
    .A2(_12480_),
    .B1(net177),
    .C1(_12492_),
    .X(_12499_));
 sky130_fd_sc_hd__a311o_4 _22545_ (.A1(_12488_),
    .A2(_12489_),
    .A3(net335),
    .B1(_12490_),
    .C1(net175),
    .X(_12500_));
 sky130_fd_sc_hd__a31o_1 _22546_ (.A1(_12057_),
    .A2(_12059_),
    .A3(_12065_),
    .B1(_12061_),
    .X(_12501_));
 sky130_fd_sc_hd__a31oi_4 _22547_ (.A1(_12057_),
    .A2(_12059_),
    .A3(_12065_),
    .B1(_12061_),
    .Y(_12502_));
 sky130_fd_sc_hd__o2111ai_4 _22548_ (.A1(_12064_),
    .A2(_12060_),
    .B1(_12062_),
    .C1(_12498_),
    .D1(_12500_),
    .Y(_12503_));
 sky130_fd_sc_hd__o21ai_2 _22549_ (.A1(_12497_),
    .A2(_12499_),
    .B1(_12501_),
    .Y(_12504_));
 sky130_fd_sc_hd__a21oi_2 _22550_ (.A1(_12491_),
    .A2(_12492_),
    .B1(net332),
    .Y(_12506_));
 sky130_fd_sc_hd__or3_1 _22551_ (.A(_11046_),
    .B(_11057_),
    .C(_12495_),
    .X(_12507_));
 sky130_fd_sc_hd__o221ai_4 _22552_ (.A1(_12064_),
    .A2(_12060_),
    .B1(_12499_),
    .B2(_12497_),
    .C1(_12062_),
    .Y(_12508_));
 sky130_fd_sc_hd__nand3_2 _22553_ (.A(_12501_),
    .B(_12500_),
    .C(_12498_),
    .Y(_12509_));
 sky130_fd_sc_hd__a31o_1 _22554_ (.A1(_12508_),
    .A2(_12509_),
    .A3(net332),
    .B1(_12506_),
    .X(_12510_));
 sky130_fd_sc_hd__a31o_2 _22555_ (.A1(_12503_),
    .A2(_12504_),
    .A3(net332),
    .B1(_12496_),
    .X(_12511_));
 sky130_fd_sc_hd__a31oi_1 _22556_ (.A1(_12508_),
    .A2(_12509_),
    .A3(net332),
    .B1(net198),
    .Y(_12512_));
 sky130_fd_sc_hd__a311oi_2 _22557_ (.A1(_12508_),
    .A2(_12509_),
    .A3(net332),
    .B1(net198),
    .C1(_12506_),
    .Y(_12513_));
 sky130_fd_sc_hd__a311o_1 _22558_ (.A1(_12508_),
    .A2(_12509_),
    .A3(net332),
    .B1(net198),
    .C1(_12506_),
    .X(_12514_));
 sky130_fd_sc_hd__a311oi_4 _22559_ (.A1(_12503_),
    .A2(_12504_),
    .A3(net332),
    .B1(net199),
    .C1(_12496_),
    .Y(_12515_));
 sky130_fd_sc_hd__a311o_1 _22560_ (.A1(_12503_),
    .A2(_12504_),
    .A3(net332),
    .B1(net199),
    .C1(_12496_),
    .X(_12517_));
 sky130_fd_sc_hd__a21oi_1 _22561_ (.A1(_12507_),
    .A2(_12512_),
    .B1(_12515_),
    .Y(_12518_));
 sky130_fd_sc_hd__and3_1 _22562_ (.A(_10634_),
    .B(_11120_),
    .C(_11122_),
    .X(_12519_));
 sky130_fd_sc_hd__nand4b_1 _22563_ (.A_N(_10644_),
    .B(_11609_),
    .C(_12519_),
    .D(_11611_),
    .Y(_12520_));
 sky130_fd_sc_hd__nand3_2 _22564_ (.A(_12083_),
    .B(_12519_),
    .C(_11612_),
    .Y(_12521_));
 sky130_fd_sc_hd__nor3b_1 _22565_ (.A(_12520_),
    .B(_12082_),
    .C_N(_12081_),
    .Y(_12522_));
 sky130_fd_sc_hd__nand3b_4 _22566_ (.A_N(_12520_),
    .B(_12083_),
    .C(_12081_),
    .Y(_12523_));
 sky130_fd_sc_hd__o211a_1 _22567_ (.A1(_12087_),
    .A2(_12082_),
    .B1(_12081_),
    .C1(_12521_),
    .X(_12524_));
 sky130_fd_sc_hd__o211ai_4 _22568_ (.A1(_12087_),
    .A2(_12082_),
    .B1(_12081_),
    .C1(_12521_),
    .Y(_12525_));
 sky130_fd_sc_hd__o211ai_2 _22569_ (.A1(_12513_),
    .A2(_12515_),
    .B1(_12523_),
    .C1(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__o21ai_1 _22570_ (.A1(_12522_),
    .A2(_12524_),
    .B1(_12518_),
    .Y(_12528_));
 sky130_fd_sc_hd__nand4_4 _22571_ (.A(_12514_),
    .B(_12517_),
    .C(_12523_),
    .D(_12525_),
    .Y(_12529_));
 sky130_fd_sc_hd__o22ai_2 _22572_ (.A1(_12513_),
    .A2(_12515_),
    .B1(_12522_),
    .B2(_12524_),
    .Y(_12530_));
 sky130_fd_sc_hd__nand3_1 _22573_ (.A(_12530_),
    .B(net311),
    .C(_12529_),
    .Y(_12531_));
 sky130_fd_sc_hd__nor2_1 _22574_ (.A(net311),
    .B(_12511_),
    .Y(_12532_));
 sky130_fd_sc_hd__a311o_4 _22575_ (.A1(_12508_),
    .A2(_12509_),
    .A3(net332),
    .B1(net311),
    .C1(_12506_),
    .X(_12533_));
 sky130_fd_sc_hd__nand3_4 _22576_ (.A(_12528_),
    .B(net311),
    .C(_12526_),
    .Y(_12534_));
 sky130_fd_sc_hd__and3_2 _22577_ (.A(_00066_),
    .B(_12533_),
    .C(_12534_),
    .X(_12535_));
 sky130_fd_sc_hd__o211ai_4 _22578_ (.A1(_14458_),
    .A2(_00000_),
    .B1(_12533_),
    .C1(_12534_),
    .Y(_12536_));
 sky130_fd_sc_hd__o211ai_4 _22579_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_12533_),
    .C1(_12534_),
    .Y(_12537_));
 sky130_fd_sc_hd__a311oi_4 _22580_ (.A1(_12530_),
    .A2(net311),
    .A3(_12529_),
    .B1(_12532_),
    .C1(_07936_),
    .Y(_12539_));
 sky130_fd_sc_hd__o211ai_4 _22581_ (.A1(net311),
    .A2(_12511_),
    .B1(_07935_),
    .C1(_12531_),
    .Y(_12540_));
 sky130_fd_sc_hd__o221a_1 _22582_ (.A1(net224),
    .A2(_11624_),
    .B1(_11630_),
    .B2(_11632_),
    .C1(_12098_),
    .X(_12541_));
 sky130_fd_sc_hd__o221ai_4 _22583_ (.A1(net224),
    .A2(_11624_),
    .B1(_11630_),
    .B2(_11632_),
    .C1(_12098_),
    .Y(_12542_));
 sky130_fd_sc_hd__o21ai_1 _22584_ (.A1(_12079_),
    .A2(_12100_),
    .B1(_12542_),
    .Y(_12543_));
 sky130_fd_sc_hd__o2bb2ai_4 _22585_ (.A1_N(_12537_),
    .A2_N(_12540_),
    .B1(_12541_),
    .B2(_12101_),
    .Y(_12544_));
 sky130_fd_sc_hd__nand4b_4 _22586_ (.A_N(_12101_),
    .B(_12537_),
    .C(_12540_),
    .D(_12542_),
    .Y(_12545_));
 sky130_fd_sc_hd__nand3_2 _22587_ (.A(_12544_),
    .B(_12545_),
    .C(net307),
    .Y(_12546_));
 sky130_fd_sc_hd__a31o_1 _22588_ (.A1(_12544_),
    .A2(_12545_),
    .A3(net307),
    .B1(_12535_),
    .X(_12547_));
 sky130_fd_sc_hd__o21bai_4 _22589_ (.A1(_12109_),
    .A2(_12115_),
    .B1_N(_12107_),
    .Y(_12548_));
 sky130_fd_sc_hd__a31o_1 _22590_ (.A1(_12544_),
    .A2(_12545_),
    .A3(net307),
    .B1(net202),
    .X(_12550_));
 sky130_fd_sc_hd__a311oi_4 _22591_ (.A1(_12544_),
    .A2(_12545_),
    .A3(net307),
    .B1(net202),
    .C1(_12535_),
    .Y(_12551_));
 sky130_fd_sc_hd__a2bb2oi_4 _22592_ (.A1_N(_07555_),
    .A2_N(_07557_),
    .B1(_12536_),
    .B2(_12546_),
    .Y(_12552_));
 sky130_fd_sc_hd__a22o_1 _22593_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_12536_),
    .B2(_12546_),
    .X(_12553_));
 sky130_fd_sc_hd__o211ai_4 _22594_ (.A1(_12535_),
    .A2(_12550_),
    .B1(_12553_),
    .C1(_12548_),
    .Y(_12554_));
 sky130_fd_sc_hd__o221ai_4 _22595_ (.A1(_12109_),
    .A2(_12115_),
    .B1(_12551_),
    .B2(_12552_),
    .C1(_12108_),
    .Y(_12555_));
 sky130_fd_sc_hd__a21oi_2 _22596_ (.A1(_12536_),
    .A2(_12546_),
    .B1(net279),
    .Y(_12556_));
 sky130_fd_sc_hd__inv_2 _22597_ (.A(_12556_),
    .Y(_12557_));
 sky130_fd_sc_hd__nand3_2 _22598_ (.A(_12554_),
    .B(_12555_),
    .C(net279),
    .Y(_12558_));
 sky130_fd_sc_hd__a31oi_4 _22599_ (.A1(_12554_),
    .A2(_12555_),
    .A3(net279),
    .B1(_12556_),
    .Y(_12559_));
 sky130_fd_sc_hd__a2bb2oi_4 _22600_ (.A1_N(_07242_),
    .A2_N(_07243_),
    .B1(_12557_),
    .B2(_12558_),
    .Y(_12561_));
 sky130_fd_sc_hd__a2bb2o_1 _22601_ (.A1_N(_07242_),
    .A2_N(_07243_),
    .B1(_12557_),
    .B2(_12558_),
    .X(_12562_));
 sky130_fd_sc_hd__o211a_2 _22602_ (.A1(_07244_),
    .A2(_07245_),
    .B1(_12557_),
    .C1(_12558_),
    .X(_12563_));
 sky130_fd_sc_hd__a311o_4 _22603_ (.A1(_12554_),
    .A2(_12555_),
    .A3(net279),
    .B1(_12556_),
    .C1(net222),
    .X(_12564_));
 sky130_fd_sc_hd__o211ai_4 _22604_ (.A1(_12137_),
    .A2(_10227_),
    .B1(_12128_),
    .C1(_12136_),
    .Y(_12565_));
 sky130_fd_sc_hd__o2111ai_4 _22605_ (.A1(_12124_),
    .A2(_12140_),
    .B1(_12562_),
    .C1(_12564_),
    .D1(_12128_),
    .Y(_12566_));
 sky130_fd_sc_hd__o211ai_4 _22606_ (.A1(_12561_),
    .A2(_12563_),
    .B1(_12125_),
    .C1(_12142_),
    .Y(_12567_));
 sky130_fd_sc_hd__nand3_2 _22607_ (.A(_12566_),
    .B(_12567_),
    .C(net277),
    .Y(_12568_));
 sky130_fd_sc_hd__a211o_2 _22608_ (.A1(_12557_),
    .A2(_12558_),
    .B1(net302),
    .C1(_04019_),
    .X(_12569_));
 sky130_fd_sc_hd__inv_2 _22609_ (.A(_12569_),
    .Y(_12570_));
 sky130_fd_sc_hd__o31a_1 _22610_ (.A1(net302),
    .A2(_04019_),
    .A3(_12559_),
    .B1(_12568_),
    .X(_12572_));
 sky130_fd_sc_hd__a31o_2 _22611_ (.A1(_12566_),
    .A2(_12567_),
    .A3(net277),
    .B1(_12570_),
    .X(_12573_));
 sky130_fd_sc_hd__a311o_1 _22612_ (.A1(_12566_),
    .A2(_12567_),
    .A3(net277),
    .B1(_12570_),
    .C1(net272),
    .X(_12574_));
 sky130_fd_sc_hd__a22oi_4 _22613_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_12568_),
    .B2(_12569_),
    .Y(_12575_));
 sky130_fd_sc_hd__a22o_2 _22614_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_12568_),
    .B2(_12569_),
    .X(_12576_));
 sky130_fd_sc_hd__a31oi_1 _22615_ (.A1(_12566_),
    .A2(_12567_),
    .A3(net277),
    .B1(net225),
    .Y(_12577_));
 sky130_fd_sc_hd__a31o_1 _22616_ (.A1(_12566_),
    .A2(_12567_),
    .A3(net277),
    .B1(net225),
    .X(_12578_));
 sky130_fd_sc_hd__and3_1 _22617_ (.A(_12568_),
    .B(_12569_),
    .C(net227),
    .X(_12579_));
 sky130_fd_sc_hd__a311o_2 _22618_ (.A1(_12566_),
    .A2(_12567_),
    .A3(net277),
    .B1(net225),
    .C1(_12570_),
    .X(_12580_));
 sky130_fd_sc_hd__a21oi_2 _22619_ (.A1(_12569_),
    .A2(_12577_),
    .B1(_12575_),
    .Y(_12581_));
 sky130_fd_sc_hd__o2111ai_2 _22620_ (.A1(_10716_),
    .A2(_10702_),
    .B1(_10715_),
    .C1(_11194_),
    .D1(_11195_),
    .Y(_12583_));
 sky130_fd_sc_hd__nor3_2 _22621_ (.A(_11687_),
    .B(_12583_),
    .C(_11689_),
    .Y(_12584_));
 sky130_fd_sc_hd__nand2_1 _22622_ (.A(_12584_),
    .B(_12153_),
    .Y(_12585_));
 sky130_fd_sc_hd__a21oi_1 _22623_ (.A1(_12584_),
    .A2(_12153_),
    .B1(_12155_),
    .Y(_12586_));
 sky130_fd_sc_hd__o211ai_4 _22624_ (.A1(_12159_),
    .A2(_12152_),
    .B1(_12156_),
    .C1(_12585_),
    .Y(_12587_));
 sky130_fd_sc_hd__and4b_1 _22625_ (.A_N(_12583_),
    .B(_11690_),
    .C(_11688_),
    .D(_10713_),
    .X(_12588_));
 sky130_fd_sc_hd__o211ai_4 _22626_ (.A1(net234),
    .A2(_12147_),
    .B1(_12584_),
    .C1(_10713_),
    .Y(_12589_));
 sky130_fd_sc_hd__nand4_4 _22627_ (.A(_12584_),
    .B(_12156_),
    .C(_12153_),
    .D(_10713_),
    .Y(_12590_));
 sky130_fd_sc_hd__a22oi_2 _22628_ (.A1(_12157_),
    .A2(_12588_),
    .B1(_12586_),
    .B2(_12161_),
    .Y(_12591_));
 sky130_fd_sc_hd__o21ai_4 _22629_ (.A1(_12152_),
    .A2(_12589_),
    .B1(_12587_),
    .Y(_12592_));
 sky130_fd_sc_hd__nand2_1 _22630_ (.A(_12592_),
    .B(_12581_),
    .Y(_12594_));
 sky130_fd_sc_hd__o221ai_2 _22631_ (.A1(_12589_),
    .A2(_12152_),
    .B1(_12575_),
    .B2(_12579_),
    .C1(_12587_),
    .Y(_12595_));
 sky130_fd_sc_hd__nand4_4 _22632_ (.A(_12576_),
    .B(_12580_),
    .C(_12587_),
    .D(_12590_),
    .Y(_12596_));
 sky130_fd_sc_hd__o21ai_1 _22633_ (.A1(_12575_),
    .A2(_12579_),
    .B1(_12592_),
    .Y(_12597_));
 sky130_fd_sc_hd__nand3_2 _22634_ (.A(_12594_),
    .B(_12595_),
    .C(net272),
    .Y(_12598_));
 sky130_fd_sc_hd__a21oi_2 _22635_ (.A1(_12568_),
    .A2(_12569_),
    .B1(net272),
    .Y(_12599_));
 sky130_fd_sc_hd__inv_2 _22636_ (.A(_12599_),
    .Y(_12600_));
 sky130_fd_sc_hd__o221ai_4 _22637_ (.A1(net296),
    .A2(_05232_),
    .B1(_12581_),
    .B2(_12591_),
    .C1(_12596_),
    .Y(_12601_));
 sky130_fd_sc_hd__and3_2 _22638_ (.A(_05486_),
    .B(_12574_),
    .C(_12598_),
    .X(_12602_));
 sky130_fd_sc_hd__a211o_2 _22639_ (.A1(_12600_),
    .A2(_12601_),
    .B1(net270),
    .C1(_05483_),
    .X(_12603_));
 sky130_fd_sc_hd__a311oi_4 _22640_ (.A1(_12597_),
    .A2(net272),
    .A3(_12596_),
    .B1(_12599_),
    .C1(net232),
    .Y(_12605_));
 sky130_fd_sc_hd__nand3_4 _22641_ (.A(_12601_),
    .B(net234),
    .C(_12600_),
    .Y(_12606_));
 sky130_fd_sc_hd__o211ai_4 _22642_ (.A1(_12573_),
    .A2(net272),
    .B1(net232),
    .C1(_12598_),
    .Y(_12607_));
 sky130_fd_sc_hd__o221a_1 _22643_ (.A1(_11707_),
    .A2(_11702_),
    .B1(_06314_),
    .B2(_12164_),
    .C1(_11701_),
    .X(_12608_));
 sky130_fd_sc_hd__a21o_1 _22644_ (.A1(_12168_),
    .A2(_12171_),
    .B1(_12172_),
    .X(_12609_));
 sky130_fd_sc_hd__a21oi_2 _22645_ (.A1(_12168_),
    .A2(_12171_),
    .B1(_12172_),
    .Y(_12610_));
 sky130_fd_sc_hd__o2bb2ai_4 _22646_ (.A1_N(_12606_),
    .A2_N(_12607_),
    .B1(_12608_),
    .B2(_12170_),
    .Y(_12611_));
 sky130_fd_sc_hd__nand3_4 _22647_ (.A(_12609_),
    .B(_12607_),
    .C(_12606_),
    .Y(_12612_));
 sky130_fd_sc_hd__nand3_1 _22648_ (.A(_12611_),
    .B(_12612_),
    .C(net245),
    .Y(_12613_));
 sky130_fd_sc_hd__a31oi_4 _22649_ (.A1(_12611_),
    .A2(_12612_),
    .A3(net245),
    .B1(_12602_),
    .Y(_12614_));
 sky130_fd_sc_hd__a31o_1 _22650_ (.A1(_12611_),
    .A2(_12612_),
    .A3(net245),
    .B1(_12602_),
    .X(_12616_));
 sky130_fd_sc_hd__o211a_1 _22651_ (.A1(_11725_),
    .A2(_11721_),
    .B1(_11719_),
    .C1(_12183_),
    .X(_12617_));
 sky130_fd_sc_hd__a22oi_2 _22652_ (.A1(_12179_),
    .A2(_12184_),
    .B1(_12190_),
    .B2(_12183_),
    .Y(_12618_));
 sky130_fd_sc_hd__a22o_1 _22653_ (.A1(_12179_),
    .A2(_12184_),
    .B1(_12190_),
    .B2(_12183_),
    .X(_12619_));
 sky130_fd_sc_hd__a31oi_2 _22654_ (.A1(_12611_),
    .A2(_12612_),
    .A3(net245),
    .B1(net252),
    .Y(_12620_));
 sky130_fd_sc_hd__a311oi_4 _22655_ (.A1(_12611_),
    .A2(_12612_),
    .A3(net245),
    .B1(net251),
    .C1(_12602_),
    .Y(_12621_));
 sky130_fd_sc_hd__a311o_1 _22656_ (.A1(_12611_),
    .A2(_12612_),
    .A3(net245),
    .B1(net252),
    .C1(_12602_),
    .X(_12622_));
 sky130_fd_sc_hd__a2bb2oi_4 _22657_ (.A1_N(net284),
    .A2_N(_06307_),
    .B1(_12603_),
    .B2(_12613_),
    .Y(_12623_));
 sky130_fd_sc_hd__a22o_1 _22658_ (.A1(_06306_),
    .A2(_06308_),
    .B1(_12603_),
    .B2(_12613_),
    .X(_12624_));
 sky130_fd_sc_hd__o211ai_1 _22659_ (.A1(_12185_),
    .A2(_12617_),
    .B1(_12622_),
    .C1(_12624_),
    .Y(_12625_));
 sky130_fd_sc_hd__o21ai_1 _22660_ (.A1(_12621_),
    .A2(_12623_),
    .B1(_12618_),
    .Y(_12627_));
 sky130_fd_sc_hd__o211ai_2 _22661_ (.A1(_05750_),
    .A2(net264),
    .B1(_12625_),
    .C1(_12627_),
    .Y(_12628_));
 sky130_fd_sc_hd__or3_1 _22662_ (.A(_05750_),
    .B(net264),
    .C(_12614_),
    .X(_12629_));
 sky130_fd_sc_hd__o21ai_1 _22663_ (.A1(_06314_),
    .A2(_12614_),
    .B1(_12618_),
    .Y(_12630_));
 sky130_fd_sc_hd__o22ai_2 _22664_ (.A1(_12185_),
    .A2(_12617_),
    .B1(_12621_),
    .B2(_12623_),
    .Y(_12631_));
 sky130_fd_sc_hd__o221ai_4 _22665_ (.A1(_05750_),
    .A2(net264),
    .B1(_12621_),
    .B2(_12630_),
    .C1(_12631_),
    .Y(_12632_));
 sky130_fd_sc_hd__o31a_1 _22666_ (.A1(_05750_),
    .A2(net264),
    .A3(_12614_),
    .B1(_12632_),
    .X(_12633_));
 sky130_fd_sc_hd__a2bb2oi_1 _22667_ (.A1_N(_06009_),
    .A2_N(net287),
    .B1(_12629_),
    .B2(_12632_),
    .Y(_12634_));
 sky130_fd_sc_hd__o211ai_4 _22668_ (.A1(_12616_),
    .A2(net242),
    .B1(net253),
    .C1(_12628_),
    .Y(_12635_));
 sky130_fd_sc_hd__o221a_2 _22669_ (.A1(_06011_),
    .A2(_06012_),
    .B1(_12614_),
    .B2(net242),
    .C1(_12632_),
    .X(_12636_));
 sky130_fd_sc_hd__o221ai_4 _22670_ (.A1(_06011_),
    .A2(_06012_),
    .B1(_12614_),
    .B2(net242),
    .C1(_12632_),
    .Y(_12638_));
 sky130_fd_sc_hd__o22ai_1 _22671_ (.A1(net263),
    .A2(_12196_),
    .B1(_12218_),
    .B2(_12211_),
    .Y(_12639_));
 sky130_fd_sc_hd__a31oi_2 _22672_ (.A1(_12203_),
    .A2(_12212_),
    .A3(_12215_),
    .B1(_12200_),
    .Y(_12640_));
 sky130_fd_sc_hd__o2bb2ai_1 _22673_ (.A1_N(_12201_),
    .A2_N(_12219_),
    .B1(_12634_),
    .B2(_12636_),
    .Y(_12641_));
 sky130_fd_sc_hd__o2111ai_4 _22674_ (.A1(net263),
    .A2(_12196_),
    .B1(_12219_),
    .C1(_12635_),
    .D1(_12638_),
    .Y(_12642_));
 sky130_fd_sc_hd__o21ai_2 _22675_ (.A1(_12634_),
    .A2(_12636_),
    .B1(_12640_),
    .Y(_12643_));
 sky130_fd_sc_hd__nand3_1 _22676_ (.A(_12639_),
    .B(_12638_),
    .C(_12635_),
    .Y(_12644_));
 sky130_fd_sc_hd__a22oi_4 _22677_ (.A1(_05991_),
    .A2(_05993_),
    .B1(_12641_),
    .B2(_12642_),
    .Y(_12645_));
 sky130_fd_sc_hd__o211ai_4 _22678_ (.A1(net260),
    .A2(net258),
    .B1(_12643_),
    .C1(_12644_),
    .Y(_12646_));
 sky130_fd_sc_hd__o211a_1 _22679_ (.A1(net242),
    .A2(_12616_),
    .B1(_05995_),
    .C1(_12628_),
    .X(_12647_));
 sky130_fd_sc_hd__or3_1 _22680_ (.A(net260),
    .B(net258),
    .C(_12633_),
    .X(_12649_));
 sky130_fd_sc_hd__o31a_1 _22681_ (.A1(net260),
    .A2(net258),
    .A3(_12633_),
    .B1(_12646_),
    .X(_12650_));
 sky130_fd_sc_hd__inv_2 _22682_ (.A(_12650_),
    .Y(_12651_));
 sky130_fd_sc_hd__a22oi_2 _22683_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_12646_),
    .B2(_12649_),
    .Y(_12652_));
 sky130_fd_sc_hd__o22ai_4 _22684_ (.A1(_05760_),
    .A2(_05762_),
    .B1(_12645_),
    .B2(_12647_),
    .Y(_12653_));
 sky130_fd_sc_hd__a31oi_1 _22685_ (.A1(net240),
    .A2(_12643_),
    .A3(_12644_),
    .B1(net261),
    .Y(_12654_));
 sky130_fd_sc_hd__o221ai_4 _22686_ (.A1(_05765_),
    .A2(_05766_),
    .B1(net240),
    .B2(_12633_),
    .C1(_12646_),
    .Y(_12655_));
 sky130_fd_sc_hd__a21oi_2 _22687_ (.A1(_12649_),
    .A2(_12654_),
    .B1(_12652_),
    .Y(_12656_));
 sky130_fd_sc_hd__nand2_1 _22688_ (.A(_12653_),
    .B(_12655_),
    .Y(_12657_));
 sky130_fd_sc_hd__and3_1 _22689_ (.A(_11273_),
    .B(_11275_),
    .C(_10798_),
    .X(_12658_));
 sky130_fd_sc_hd__nand3_1 _22690_ (.A(_12228_),
    .B(_12658_),
    .C(_11766_),
    .Y(_12660_));
 sky130_fd_sc_hd__o211ai_4 _22691_ (.A1(_12233_),
    .A2(_12227_),
    .B1(_12230_),
    .C1(_12660_),
    .Y(_12661_));
 sky130_fd_sc_hd__and4b_1 _22692_ (.A_N(_10795_),
    .B(_11763_),
    .C(_12658_),
    .D(_11765_),
    .X(_12662_));
 sky130_fd_sc_hd__nand3_4 _22693_ (.A(_12662_),
    .B(_12230_),
    .C(_12228_),
    .Y(_12663_));
 sky130_fd_sc_hd__nand2_1 _22694_ (.A(_12661_),
    .B(_12663_),
    .Y(_12664_));
 sky130_fd_sc_hd__a21oi_2 _22695_ (.A1(_12661_),
    .A2(_12663_),
    .B1(_12657_),
    .Y(_12665_));
 sky130_fd_sc_hd__o22ai_4 _22696_ (.A1(_06291_),
    .A2(_06292_),
    .B1(_12656_),
    .B2(_12664_),
    .Y(_12666_));
 sky130_fd_sc_hd__o22a_1 _22697_ (.A1(_06286_),
    .A2(_06288_),
    .B1(_12645_),
    .B2(_12647_),
    .X(_12667_));
 sky130_fd_sc_hd__or3_1 _22698_ (.A(_06291_),
    .B(_06292_),
    .C(_12650_),
    .X(_12668_));
 sky130_fd_sc_hd__a22o_1 _22699_ (.A1(_12653_),
    .A2(_12655_),
    .B1(_12661_),
    .B2(_12663_),
    .X(_12669_));
 sky130_fd_sc_hd__nand3_2 _22700_ (.A(_12655_),
    .B(_12661_),
    .C(_12663_),
    .Y(_12671_));
 sky130_fd_sc_hd__nand4_2 _22701_ (.A(_12653_),
    .B(_12655_),
    .C(_12661_),
    .D(_12663_),
    .Y(_12672_));
 sky130_fd_sc_hd__nand3_2 _22702_ (.A(_12669_),
    .B(_12672_),
    .C(net213),
    .Y(_12673_));
 sky130_fd_sc_hd__a311oi_4 _22703_ (.A1(_12669_),
    .A2(_12672_),
    .A3(net213),
    .B1(_12667_),
    .C1(net292),
    .Y(_12674_));
 sky130_fd_sc_hd__nand3_4 _22704_ (.A(_12673_),
    .B(_05507_),
    .C(_12668_),
    .Y(_12675_));
 sky130_fd_sc_hd__o221ai_4 _22705_ (.A1(net213),
    .A2(_12651_),
    .B1(_12665_),
    .B2(_12666_),
    .C1(net292),
    .Y(_12676_));
 sky130_fd_sc_hd__o22a_1 _22706_ (.A1(net295),
    .A2(_12238_),
    .B1(_12240_),
    .B2(_11779_),
    .X(_12677_));
 sky130_fd_sc_hd__a21o_1 _22707_ (.A1(_12245_),
    .A2(_12243_),
    .B1(_12246_),
    .X(_12678_));
 sky130_fd_sc_hd__a21oi_1 _22708_ (.A1(_12245_),
    .A2(_12243_),
    .B1(_12246_),
    .Y(_12679_));
 sky130_fd_sc_hd__o2bb2ai_4 _22709_ (.A1_N(_12675_),
    .A2_N(_12676_),
    .B1(_12677_),
    .B2(_12244_),
    .Y(_12680_));
 sky130_fd_sc_hd__nand3_4 _22710_ (.A(_12678_),
    .B(_12676_),
    .C(_12675_),
    .Y(_12682_));
 sky130_fd_sc_hd__nand3_1 _22711_ (.A(_12680_),
    .B(_12682_),
    .C(net210),
    .Y(_12683_));
 sky130_fd_sc_hd__o221a_4 _22712_ (.A1(net213),
    .A2(_12651_),
    .B1(_12665_),
    .B2(_12666_),
    .C1(_06613_),
    .X(_12684_));
 sky130_fd_sc_hd__a211o_1 _22713_ (.A1(_12668_),
    .A2(_12673_),
    .B1(_06608_),
    .C1(_06610_),
    .X(_12685_));
 sky130_fd_sc_hd__a31oi_4 _22714_ (.A1(_12680_),
    .A2(_12682_),
    .A3(net210),
    .B1(_12684_),
    .Y(_12686_));
 sky130_fd_sc_hd__inv_2 _22715_ (.A(_12686_),
    .Y(_12687_));
 sky130_fd_sc_hd__a31oi_2 _22716_ (.A1(_04238_),
    .A2(_12239_),
    .A3(_12251_),
    .B1(_12263_),
    .Y(_12688_));
 sky130_fd_sc_hd__o21a_1 _22717_ (.A1(_11791_),
    .A2(_11806_),
    .B1(_12261_),
    .X(_12689_));
 sky130_fd_sc_hd__o21ai_2 _22718_ (.A1(_11791_),
    .A2(_11806_),
    .B1(_12261_),
    .Y(_12690_));
 sky130_fd_sc_hd__o21ai_1 _22719_ (.A1(net299),
    .A2(_12257_),
    .B1(_12690_),
    .Y(_12691_));
 sky130_fd_sc_hd__a31o_1 _22720_ (.A1(_12680_),
    .A2(_12682_),
    .A3(net210),
    .B1(net294),
    .X(_12693_));
 sky130_fd_sc_hd__a311oi_4 _22721_ (.A1(_12680_),
    .A2(_12682_),
    .A3(net210),
    .B1(_12684_),
    .C1(net294),
    .Y(_12694_));
 sky130_fd_sc_hd__a22oi_4 _22722_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_12683_),
    .B2(_12685_),
    .Y(_12695_));
 sky130_fd_sc_hd__a22o_1 _22723_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_12683_),
    .B2(_12685_),
    .X(_12696_));
 sky130_fd_sc_hd__o221ai_1 _22724_ (.A1(_12260_),
    .A2(_12688_),
    .B1(_12693_),
    .B2(_12684_),
    .C1(_12696_),
    .Y(_12697_));
 sky130_fd_sc_hd__o22ai_1 _22725_ (.A1(_12258_),
    .A2(_12689_),
    .B1(_12694_),
    .B2(_12695_),
    .Y(_12698_));
 sky130_fd_sc_hd__nand3_1 _22726_ (.A(_12697_),
    .B(_12698_),
    .C(net208),
    .Y(_12699_));
 sky130_fd_sc_hd__or3_1 _22727_ (.A(net230),
    .B(_06901_),
    .C(_12686_),
    .X(_12700_));
 sky130_fd_sc_hd__o21ai_1 _22728_ (.A1(net295),
    .A2(_12686_),
    .B1(_12691_),
    .Y(_12701_));
 sky130_fd_sc_hd__o22ai_2 _22729_ (.A1(_12260_),
    .A2(_12688_),
    .B1(_12694_),
    .B2(_12695_),
    .Y(_12702_));
 sky130_fd_sc_hd__o221ai_4 _22730_ (.A1(_06899_),
    .A2(_06901_),
    .B1(_12694_),
    .B2(_12701_),
    .C1(_12702_),
    .Y(_12704_));
 sky130_fd_sc_hd__o31a_2 _22731_ (.A1(net230),
    .A2(_06901_),
    .A3(_12686_),
    .B1(_12704_),
    .X(_12705_));
 sky130_fd_sc_hd__inv_2 _22732_ (.A(_12705_),
    .Y(_12706_));
 sky130_fd_sc_hd__o211ai_4 _22733_ (.A1(_12687_),
    .A2(net208),
    .B1(_04238_),
    .C1(_12699_),
    .Y(_12707_));
 sky130_fd_sc_hd__o211a_2 _22734_ (.A1(net208),
    .A2(_12686_),
    .B1(net299),
    .C1(_12704_),
    .X(_12708_));
 sky130_fd_sc_hd__nand3_2 _22735_ (.A(_12704_),
    .B(net299),
    .C(_12700_),
    .Y(_12709_));
 sky130_fd_sc_hd__nand2_1 _22736_ (.A(_12707_),
    .B(_12709_),
    .Y(_12710_));
 sky130_fd_sc_hd__o2bb2ai_2 _22737_ (.A1_N(_11957_),
    .A2_N(_11958_),
    .B1(_12271_),
    .B2(_02137_),
    .Y(_12711_));
 sky130_fd_sc_hd__a31oi_4 _22738_ (.A1(_11957_),
    .A2(_11958_),
    .A3(_12277_),
    .B1(_12273_),
    .Y(_12712_));
 sky130_fd_sc_hd__a22oi_4 _22739_ (.A1(_12707_),
    .A2(_12709_),
    .B1(_12711_),
    .B2(_12277_),
    .Y(_12713_));
 sky130_fd_sc_hd__o2111a_1 _22740_ (.A1(_02148_),
    .A2(_12272_),
    .B1(_12707_),
    .C1(_12709_),
    .D1(_12711_),
    .X(_12715_));
 sky130_fd_sc_hd__o22ai_4 _22741_ (.A1(_07227_),
    .A2(_07229_),
    .B1(_12713_),
    .B2(_12715_),
    .Y(_12716_));
 sky130_fd_sc_hd__o21ai_4 _22742_ (.A1(_12712_),
    .A2(_12710_),
    .B1(net185),
    .Y(_12717_));
 sky130_fd_sc_hd__o22ai_4 _22743_ (.A1(net185),
    .A2(_12705_),
    .B1(_12713_),
    .B2(_12717_),
    .Y(_12718_));
 sky130_fd_sc_hd__o22a_1 _22744_ (.A1(net185),
    .A2(_12705_),
    .B1(_12713_),
    .B2(_12717_),
    .X(_12719_));
 sky130_fd_sc_hd__o311a_1 _22745_ (.A1(_07227_),
    .A2(_07229_),
    .A3(_12706_),
    .B1(_12716_),
    .C1(_02148_),
    .X(_12720_));
 sky130_fd_sc_hd__o211ai_4 _22746_ (.A1(_12706_),
    .A2(net185),
    .B1(_02148_),
    .C1(_12716_),
    .Y(_12721_));
 sky130_fd_sc_hd__o221a_1 _22747_ (.A1(net185),
    .A2(_12705_),
    .B1(_12713_),
    .B2(_12717_),
    .C1(_02137_),
    .X(_12722_));
 sky130_fd_sc_hd__o221ai_4 _22748_ (.A1(net185),
    .A2(_12705_),
    .B1(_12713_),
    .B2(_12717_),
    .C1(_02137_),
    .Y(_12723_));
 sky130_fd_sc_hd__and4_1 _22749_ (.A(_10851_),
    .B(_10852_),
    .C(_11347_),
    .D(_11348_),
    .X(_12724_));
 sky130_fd_sc_hd__nand3_1 _22750_ (.A(_12292_),
    .B(_12724_),
    .C(_11837_),
    .Y(_12726_));
 sky130_fd_sc_hd__o211ai_4 _22751_ (.A1(_12296_),
    .A2(_12291_),
    .B1(_12294_),
    .C1(_12726_),
    .Y(_12727_));
 sky130_fd_sc_hd__nor4b_1 _22752_ (.A(_10855_),
    .B(_11832_),
    .C(_11834_),
    .D_N(_12724_),
    .Y(_12728_));
 sky130_fd_sc_hd__nand3_4 _22753_ (.A(_12728_),
    .B(_12294_),
    .C(_12292_),
    .Y(_12729_));
 sky130_fd_sc_hd__nand2_2 _22754_ (.A(_12727_),
    .B(_12729_),
    .Y(_12730_));
 sky130_fd_sc_hd__inv_2 _22755_ (.A(_12730_),
    .Y(_12731_));
 sky130_fd_sc_hd__a22o_2 _22756_ (.A1(_12721_),
    .A2(_12723_),
    .B1(_12727_),
    .B2(_12729_),
    .X(_12732_));
 sky130_fd_sc_hd__o211a_1 _22757_ (.A1(_12718_),
    .A2(_02148_),
    .B1(_12729_),
    .C1(_12727_),
    .X(_12733_));
 sky130_fd_sc_hd__o2111ai_4 _22758_ (.A1(_02148_),
    .A2(_12718_),
    .B1(_12721_),
    .C1(_12727_),
    .D1(_12729_),
    .Y(_12734_));
 sky130_fd_sc_hd__nand3_1 _22759_ (.A(_12732_),
    .B(_12734_),
    .C(net163),
    .Y(_12735_));
 sky130_fd_sc_hd__o311a_2 _22760_ (.A1(_07227_),
    .A2(_07229_),
    .A3(_12706_),
    .B1(_12716_),
    .C1(_07550_),
    .X(_12736_));
 sky130_fd_sc_hd__or3_1 _22761_ (.A(_07544_),
    .B(net184),
    .C(_12719_),
    .X(_12737_));
 sky130_fd_sc_hd__a31oi_4 _22762_ (.A1(_12732_),
    .A2(_12734_),
    .A3(net163),
    .B1(_12736_),
    .Y(_12738_));
 sky130_fd_sc_hd__a21oi_1 _22763_ (.A1(_12735_),
    .A2(_12737_),
    .B1(net161),
    .Y(_12739_));
 sky130_fd_sc_hd__or3_2 _22764_ (.A(_07912_),
    .B(_07914_),
    .C(_12738_),
    .X(_12740_));
 sky130_fd_sc_hd__a31o_1 _22765_ (.A1(_12732_),
    .A2(_12734_),
    .A3(net163),
    .B1(_00251_),
    .X(_12741_));
 sky130_fd_sc_hd__a311oi_4 _22766_ (.A1(_12732_),
    .A2(_12734_),
    .A3(net163),
    .B1(_12736_),
    .C1(_00251_),
    .Y(_12742_));
 sky130_fd_sc_hd__a31o_1 _22767_ (.A1(_07545_),
    .A2(_07547_),
    .A3(_12718_),
    .B1(_12741_),
    .X(_12743_));
 sky130_fd_sc_hd__a22oi_2 _22768_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_12735_),
    .B2(_12737_),
    .Y(_12744_));
 sky130_fd_sc_hd__a22o_1 _22769_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_12735_),
    .B2(_12737_),
    .X(_12745_));
 sky130_fd_sc_hd__a21o_1 _22770_ (.A1(_12306_),
    .A2(_12309_),
    .B1(_12310_),
    .X(_12747_));
 sky130_fd_sc_hd__a21oi_2 _22771_ (.A1(_12306_),
    .A2(_12309_),
    .B1(_12310_),
    .Y(_12748_));
 sky130_fd_sc_hd__o21a_1 _22772_ (.A1(_12742_),
    .A2(_12744_),
    .B1(_12748_),
    .X(_12749_));
 sky130_fd_sc_hd__o21ai_2 _22773_ (.A1(_12742_),
    .A2(_12744_),
    .B1(_12748_),
    .Y(_12750_));
 sky130_fd_sc_hd__o21ai_2 _22774_ (.A1(_00240_),
    .A2(_12738_),
    .B1(_12747_),
    .Y(_12751_));
 sky130_fd_sc_hd__o211ai_2 _22775_ (.A1(_12736_),
    .A2(_12741_),
    .B1(_12747_),
    .C1(_12745_),
    .Y(_12752_));
 sky130_fd_sc_hd__o22ai_4 _22776_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_12742_),
    .B2(_12751_),
    .Y(_12753_));
 sky130_fd_sc_hd__o211ai_4 _22777_ (.A1(_12742_),
    .A2(_12751_),
    .B1(net161),
    .C1(_12750_),
    .Y(_12754_));
 sky130_fd_sc_hd__o22a_1 _22778_ (.A1(net161),
    .A2(_12738_),
    .B1(_12749_),
    .B2(_12753_),
    .X(_12755_));
 sky130_fd_sc_hd__o22ai_4 _22779_ (.A1(net161),
    .A2(_12738_),
    .B1(_12749_),
    .B2(_12753_),
    .Y(_12756_));
 sky130_fd_sc_hd__o221a_2 _22780_ (.A1(_11861_),
    .A2(_11864_),
    .B1(_11298_),
    .B2(_12322_),
    .C1(_11860_),
    .X(_12758_));
 sky130_fd_sc_hd__o311a_1 _22781_ (.A1(_11383_),
    .A2(_11859_),
    .A3(_11863_),
    .B1(_12326_),
    .C1(_11862_),
    .X(_12759_));
 sky130_fd_sc_hd__a21o_1 _22782_ (.A1(_12326_),
    .A2(_12328_),
    .B1(_12323_),
    .X(_12760_));
 sky130_fd_sc_hd__o22a_1 _22783_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_12749_),
    .B2(_12753_),
    .X(_12761_));
 sky130_fd_sc_hd__a311oi_4 _22784_ (.A1(_12750_),
    .A2(_12752_),
    .A3(net161),
    .B1(_12739_),
    .C1(_12899_),
    .Y(_12762_));
 sky130_fd_sc_hd__o221ai_4 _22785_ (.A1(_12867_),
    .A2(_12877_),
    .B1(net161),
    .B2(_12738_),
    .C1(_12754_),
    .Y(_12763_));
 sky130_fd_sc_hd__a2bb2oi_4 _22786_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_12740_),
    .B2(_12754_),
    .Y(_12764_));
 sky130_fd_sc_hd__o21ai_2 _22787_ (.A1(net361),
    .A2(net345),
    .B1(_12756_),
    .Y(_12765_));
 sky130_fd_sc_hd__o211ai_1 _22788_ (.A1(_12325_),
    .A2(_12758_),
    .B1(_12763_),
    .C1(_12765_),
    .Y(_12766_));
 sky130_fd_sc_hd__o22ai_1 _22789_ (.A1(_12323_),
    .A2(_12759_),
    .B1(_12762_),
    .B2(_12764_),
    .Y(_12767_));
 sky130_fd_sc_hd__o211ai_2 _22790_ (.A1(net180),
    .A2(_08298_),
    .B1(_12766_),
    .C1(_12767_),
    .Y(_12769_));
 sky130_fd_sc_hd__and3_1 _22791_ (.A(_08297_),
    .B(_08299_),
    .C(_12756_),
    .X(_12770_));
 sky130_fd_sc_hd__or3_1 _22792_ (.A(net180),
    .B(_08298_),
    .C(_12755_),
    .X(_12771_));
 sky130_fd_sc_hd__nand3_2 _22793_ (.A(_12765_),
    .B(_12760_),
    .C(_12763_),
    .Y(_12772_));
 sky130_fd_sc_hd__o22ai_4 _22794_ (.A1(_12325_),
    .A2(_12758_),
    .B1(_12762_),
    .B2(_12764_),
    .Y(_12773_));
 sky130_fd_sc_hd__nand3_2 _22795_ (.A(_12773_),
    .B(_08300_),
    .C(_12772_),
    .Y(_12774_));
 sky130_fd_sc_hd__o21ai_1 _22796_ (.A1(_08300_),
    .A2(_12755_),
    .B1(_12774_),
    .Y(_12775_));
 sky130_fd_sc_hd__a31oi_4 _22797_ (.A1(_12773_),
    .A2(_08300_),
    .A3(_12772_),
    .B1(_12770_),
    .Y(_12776_));
 sky130_fd_sc_hd__o221a_2 _22798_ (.A1(_08705_),
    .A2(_08707_),
    .B1(_12755_),
    .B2(_08300_),
    .C1(_12774_),
    .X(_12777_));
 sky130_fd_sc_hd__o211a_1 _22799_ (.A1(_12756_),
    .A2(_08300_),
    .B1(_11309_),
    .C1(_12769_),
    .X(_12778_));
 sky130_fd_sc_hd__o211ai_4 _22800_ (.A1(_12756_),
    .A2(_08300_),
    .B1(_11309_),
    .C1(_12769_),
    .Y(_12780_));
 sky130_fd_sc_hd__and3_1 _22801_ (.A(_12771_),
    .B(_12774_),
    .C(_11298_),
    .X(_12781_));
 sky130_fd_sc_hd__o211ai_2 _22802_ (.A1(_08300_),
    .A2(_12755_),
    .B1(_11298_),
    .C1(_12774_),
    .Y(_12782_));
 sky130_fd_sc_hd__o311a_1 _22803_ (.A1(_11399_),
    .A2(_11876_),
    .A3(_11878_),
    .B1(_11882_),
    .C1(_12340_),
    .X(_12783_));
 sky130_fd_sc_hd__o21ai_2 _22804_ (.A1(_11951_),
    .A2(_12339_),
    .B1(_12344_),
    .Y(_12784_));
 sky130_fd_sc_hd__a32o_1 _22805_ (.A1(_09982_),
    .A2(_10004_),
    .A3(_12338_),
    .B1(_12344_),
    .B2(_11951_),
    .X(_12785_));
 sky130_fd_sc_hd__o2bb2ai_1 _22806_ (.A1_N(_12780_),
    .A2_N(_12782_),
    .B1(_12783_),
    .B2(_12343_),
    .Y(_12786_));
 sky130_fd_sc_hd__o2111ai_4 _22807_ (.A1(_11951_),
    .A2(_12339_),
    .B1(_12344_),
    .C1(_12780_),
    .D1(_12782_),
    .Y(_12787_));
 sky130_fd_sc_hd__a21oi_2 _22808_ (.A1(_12786_),
    .A2(_12787_),
    .B1(_08715_),
    .Y(_12788_));
 sky130_fd_sc_hd__or3_1 _22809_ (.A(net158),
    .B(_08712_),
    .C(_12776_),
    .X(_12789_));
 sky130_fd_sc_hd__nand3_2 _22810_ (.A(_12786_),
    .B(_12787_),
    .C(_08714_),
    .Y(_12791_));
 sky130_fd_sc_hd__a2bb2oi_2 _22811_ (.A1_N(_09927_),
    .A2_N(_09949_),
    .B1(_12789_),
    .B2(_12791_),
    .Y(_12792_));
 sky130_fd_sc_hd__a22o_1 _22812_ (.A1(_09938_),
    .A2(_09960_),
    .B1(_12789_),
    .B2(_12791_),
    .X(_12793_));
 sky130_fd_sc_hd__o221a_1 _22813_ (.A1(net365),
    .A2(net362),
    .B1(_08714_),
    .B2(_12776_),
    .C1(_12791_),
    .X(_12794_));
 sky130_fd_sc_hd__o221ai_2 _22814_ (.A1(net365),
    .A2(net362),
    .B1(_08714_),
    .B2(_12776_),
    .C1(_12791_),
    .Y(_12795_));
 sky130_fd_sc_hd__a32o_1 _22815_ (.A1(_08907_),
    .A2(_12349_),
    .A3(_12350_),
    .B1(_11892_),
    .B2(_11898_),
    .X(_12796_));
 sky130_fd_sc_hd__a21oi_2 _22816_ (.A1(_12354_),
    .A2(_12356_),
    .B1(_12357_),
    .Y(_12797_));
 sky130_fd_sc_hd__o21ai_2 _22817_ (.A1(_12353_),
    .A2(_12355_),
    .B1(_12358_),
    .Y(_12798_));
 sky130_fd_sc_hd__o21ai_1 _22818_ (.A1(_12792_),
    .A2(_12794_),
    .B1(_12797_),
    .Y(_12799_));
 sky130_fd_sc_hd__a32oi_1 _22819_ (.A1(_10015_),
    .A2(_12789_),
    .A3(_12791_),
    .B1(_12796_),
    .B2(_12358_),
    .Y(_12800_));
 sky130_fd_sc_hd__nand2_1 _22820_ (.A(_12795_),
    .B(_12798_),
    .Y(_12802_));
 sky130_fd_sc_hd__o221ai_4 _22821_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_12792_),
    .B2(_12802_),
    .C1(_12799_),
    .Y(_12803_));
 sky130_fd_sc_hd__or4_4 _22822_ (.A(_09120_),
    .B(_09121_),
    .C(_12777_),
    .D(_12788_),
    .X(_12804_));
 sky130_fd_sc_hd__o31a_2 _22823_ (.A1(_09125_),
    .A2(_12777_),
    .A3(_12788_),
    .B1(_12803_),
    .X(_12805_));
 sky130_fd_sc_hd__o21ai_2 _22824_ (.A1(_09559_),
    .A2(_09560_),
    .B1(_12805_),
    .Y(_12806_));
 sky130_fd_sc_hd__a21oi_2 _22825_ (.A1(_12370_),
    .A2(_12373_),
    .B1(_12368_),
    .Y(_12807_));
 sky130_fd_sc_hd__a21o_1 _22826_ (.A1(_12370_),
    .A2(_12373_),
    .B1(_12368_),
    .X(_12808_));
 sky130_fd_sc_hd__o311a_2 _22827_ (.A1(_09125_),
    .A2(_12777_),
    .A3(_12788_),
    .B1(_08907_),
    .C1(_12803_),
    .X(_12809_));
 sky130_fd_sc_hd__o211ai_4 _22828_ (.A1(_08863_),
    .A2(_08885_),
    .B1(_12803_),
    .C1(_12804_),
    .Y(_12810_));
 sky130_fd_sc_hd__a21oi_2 _22829_ (.A1(_12803_),
    .A2(_12804_),
    .B1(_08907_),
    .Y(_12811_));
 sky130_fd_sc_hd__a22o_1 _22830_ (.A1(_08830_),
    .A2(_08852_),
    .B1(_12803_),
    .B2(_12804_),
    .X(_12813_));
 sky130_fd_sc_hd__o211ai_2 _22831_ (.A1(_12368_),
    .A2(_12380_),
    .B1(_12810_),
    .C1(_12813_),
    .Y(_12814_));
 sky130_fd_sc_hd__o21ai_1 _22832_ (.A1(_12809_),
    .A2(_12811_),
    .B1(_12807_),
    .Y(_12815_));
 sky130_fd_sc_hd__nand3_1 _22833_ (.A(_12813_),
    .B(_12807_),
    .C(_12810_),
    .Y(_12816_));
 sky130_fd_sc_hd__o22ai_2 _22834_ (.A1(_12368_),
    .A2(_12380_),
    .B1(_12809_),
    .B2(_12811_),
    .Y(_12817_));
 sky130_fd_sc_hd__o2111ai_4 _22835_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .C1(_12816_),
    .D1(_12817_),
    .Y(_12818_));
 sky130_fd_sc_hd__or3_1 _22836_ (.A(_09553_),
    .B(net155),
    .C(_12805_),
    .X(_12819_));
 sky130_fd_sc_hd__o2111ai_4 _22837_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .C1(_12814_),
    .D1(_12815_),
    .Y(_12820_));
 sky130_fd_sc_hd__o31a_1 _22838_ (.A1(_09553_),
    .A2(net155),
    .A3(_12805_),
    .B1(_12820_),
    .X(_12821_));
 sky130_fd_sc_hd__inv_2 _22839_ (.A(_12821_),
    .Y(_12822_));
 sky130_fd_sc_hd__and3_1 _22840_ (.A(_07899_),
    .B(_12806_),
    .C(_12818_),
    .X(_12824_));
 sky130_fd_sc_hd__nand3_1 _22841_ (.A(_07899_),
    .B(_12806_),
    .C(_12818_),
    .Y(_12825_));
 sky130_fd_sc_hd__o221ai_4 _22842_ (.A1(net368),
    .A2(_07866_),
    .B1(net143),
    .B2(_12805_),
    .C1(_12820_),
    .Y(_12826_));
 sky130_fd_sc_hd__o31a_1 _22843_ (.A1(_06945_),
    .A2(_06967_),
    .A3(_12383_),
    .B1(_12386_),
    .X(_12827_));
 sky130_fd_sc_hd__o21ai_2 _22844_ (.A1(_12384_),
    .A2(_12387_),
    .B1(_12390_),
    .Y(_12828_));
 sky130_fd_sc_hd__a21oi_1 _22845_ (.A1(_12386_),
    .A2(_12388_),
    .B1(_12389_),
    .Y(_12829_));
 sky130_fd_sc_hd__o2111ai_1 _22846_ (.A1(_12384_),
    .A2(_12387_),
    .B1(_12390_),
    .C1(_12825_),
    .D1(_12826_),
    .Y(_12830_));
 sky130_fd_sc_hd__o2bb2ai_1 _22847_ (.A1_N(_12825_),
    .A2_N(_12826_),
    .B1(_12827_),
    .B2(_12389_),
    .Y(_12831_));
 sky130_fd_sc_hd__o211ai_2 _22848_ (.A1(_09571_),
    .A2(_09573_),
    .B1(_12830_),
    .C1(_12831_),
    .Y(_12832_));
 sky130_fd_sc_hd__a21o_1 _22849_ (.A1(_12825_),
    .A2(_12826_),
    .B1(_12828_),
    .X(_12833_));
 sky130_fd_sc_hd__a31oi_1 _22850_ (.A1(_07888_),
    .A2(_12819_),
    .A3(_12820_),
    .B1(_12829_),
    .Y(_12835_));
 sky130_fd_sc_hd__a31o_1 _22851_ (.A1(_07888_),
    .A2(_12819_),
    .A3(_12820_),
    .B1(_12829_),
    .X(_12836_));
 sky130_fd_sc_hd__o2111ai_4 _22852_ (.A1(_12824_),
    .A2(_12836_),
    .B1(_12833_),
    .C1(_09575_),
    .D1(_09577_),
    .Y(_12837_));
 sky130_fd_sc_hd__o21a_2 _22853_ (.A1(_09579_),
    .A2(_12822_),
    .B1(_12832_),
    .X(_12838_));
 sky130_fd_sc_hd__nand2_1 _22854_ (.A(_12395_),
    .B(_12400_),
    .Y(_12839_));
 sky130_fd_sc_hd__o221ai_4 _22855_ (.A1(_06989_),
    .A2(net375),
    .B1(_09579_),
    .B2(_12821_),
    .C1(_12837_),
    .Y(_12840_));
 sky130_fd_sc_hd__o2111ai_4 _22856_ (.A1(_12822_),
    .A2(_09579_),
    .B1(_07022_),
    .C1(net376),
    .D1(_12832_),
    .Y(_12841_));
 sky130_fd_sc_hd__a22oi_4 _22857_ (.A1(_12395_),
    .A2(_12400_),
    .B1(_12840_),
    .B2(_12841_),
    .Y(_12842_));
 sky130_fd_sc_hd__a41o_2 _22858_ (.A1(_12395_),
    .A2(_12400_),
    .A3(_12840_),
    .A4(_12841_),
    .B1(_10479_),
    .X(_12843_));
 sky130_fd_sc_hd__o21ai_1 _22859_ (.A1(_10477_),
    .A2(_10478_),
    .B1(_12838_),
    .Y(_12844_));
 sky130_fd_sc_hd__nand3_1 _22860_ (.A(_12839_),
    .B(_12840_),
    .C(_12841_),
    .Y(_12846_));
 sky130_fd_sc_hd__a21o_1 _22861_ (.A1(_12840_),
    .A2(_12841_),
    .B1(_12839_),
    .X(_12847_));
 sky130_fd_sc_hd__o211ai_1 _22862_ (.A1(_10474_),
    .A2(net138),
    .B1(_12846_),
    .C1(_12847_),
    .Y(_12848_));
 sky130_fd_sc_hd__o22ai_4 _22863_ (.A1(_10480_),
    .A2(_12838_),
    .B1(_12842_),
    .B2(_12843_),
    .Y(_12849_));
 sky130_fd_sc_hd__o221a_1 _22864_ (.A1(_10480_),
    .A2(_12838_),
    .B1(_12842_),
    .B2(_12843_),
    .C1(_06343_),
    .X(_12850_));
 sky130_fd_sc_hd__o221ai_4 _22865_ (.A1(_10480_),
    .A2(_12838_),
    .B1(_12842_),
    .B2(_12843_),
    .C1(_06343_),
    .Y(_12851_));
 sky130_fd_sc_hd__o211ai_1 _22866_ (.A1(net381),
    .A2(_06310_),
    .B1(_12844_),
    .C1(_12848_),
    .Y(_12852_));
 sky130_fd_sc_hd__o211ai_1 _22867_ (.A1(_05851_),
    .A2(_12403_),
    .B1(_12402_),
    .C1(_12401_),
    .Y(_12853_));
 sky130_fd_sc_hd__nand2_1 _22868_ (.A(_12404_),
    .B(_12853_),
    .Y(_12854_));
 sky130_fd_sc_hd__a22oi_1 _22869_ (.A1(_12851_),
    .A2(_12852_),
    .B1(_12853_),
    .B2(_12404_),
    .Y(_12855_));
 sky130_fd_sc_hd__a21oi_1 _22870_ (.A1(_12849_),
    .A2(_06332_),
    .B1(_12854_),
    .Y(_12857_));
 sky130_fd_sc_hd__a31o_1 _22871_ (.A1(_06332_),
    .A2(_12844_),
    .A3(_12848_),
    .B1(_12854_),
    .X(_12858_));
 sky130_fd_sc_hd__a211o_1 _22872_ (.A1(_12857_),
    .A2(_12851_),
    .B1(_10953_),
    .C1(_12855_),
    .X(_12859_));
 sky130_fd_sc_hd__or3_1 _22873_ (.A(_10949_),
    .B(net136),
    .C(_12849_),
    .X(_12860_));
 sky130_fd_sc_hd__a32o_1 _22874_ (.A1(_05512_),
    .A2(net396),
    .A3(_12409_),
    .B1(_12411_),
    .B2(_12408_),
    .X(_12861_));
 sky130_fd_sc_hd__a21oi_1 _22875_ (.A1(net406),
    .A2(_05840_),
    .B1(_12861_),
    .Y(_12862_));
 sky130_fd_sc_hd__o21ai_1 _22876_ (.A1(_05763_),
    .A2(_05785_),
    .B1(_12861_),
    .Y(_12863_));
 sky130_fd_sc_hd__a31o_1 _22877_ (.A1(net406),
    .A2(_05840_),
    .A3(_12861_),
    .B1(_11464_),
    .X(_12864_));
 sky130_fd_sc_hd__a211o_1 _22878_ (.A1(_12859_),
    .A2(_12860_),
    .B1(_12862_),
    .C1(_12864_),
    .X(_12865_));
 sky130_fd_sc_hd__o221ai_2 _22879_ (.A1(_10954_),
    .A2(_12849_),
    .B1(_12862_),
    .B2(_12864_),
    .C1(_12859_),
    .Y(_12866_));
 sky130_fd_sc_hd__nand2_1 _22880_ (.A(_12865_),
    .B(_12866_),
    .Y(_12868_));
 sky130_fd_sc_hd__or4_1 _22881_ (.A(_03289_),
    .B(net407),
    .C(_05218_),
    .D(_11942_),
    .X(_12869_));
 sky130_fd_sc_hd__o21ai_1 _22882_ (.A1(_12414_),
    .A2(_12415_),
    .B1(_12869_),
    .Y(_12870_));
 sky130_fd_sc_hd__o211a_1 _22883_ (.A1(_12414_),
    .A2(_12415_),
    .B1(_05545_),
    .C1(_12869_),
    .X(_12871_));
 sky130_fd_sc_hd__a21o_1 _22884_ (.A1(_12865_),
    .A2(_12866_),
    .B1(_05556_),
    .X(_12872_));
 sky130_fd_sc_hd__and3_1 _22885_ (.A(_05556_),
    .B(_12865_),
    .C(_12866_),
    .X(_12873_));
 sky130_fd_sc_hd__o21a_1 _22886_ (.A1(_11944_),
    .A2(_12871_),
    .B1(_12868_),
    .X(_12874_));
 sky130_fd_sc_hd__or3_1 _22887_ (.A(_05051_),
    .B(_12418_),
    .C(_12874_),
    .X(_12875_));
 sky130_fd_sc_hd__o21ai_1 _22888_ (.A1(_05051_),
    .A2(_12418_),
    .B1(_12874_),
    .Y(_12876_));
 sky130_fd_sc_hd__and2_1 _22889_ (.A(_12875_),
    .B(_12876_),
    .X(net91));
 sky130_fd_sc_hd__o2bb2a_1 _22890_ (.A1_N(_12418_),
    .A2_N(_12874_),
    .B1(_04832_),
    .B2(_04942_),
    .X(_12878_));
 sky130_fd_sc_hd__a32oi_4 _22891_ (.A1(_07899_),
    .A2(_12806_),
    .A3(_12818_),
    .B1(_12826_),
    .B2(_12828_),
    .Y(_12879_));
 sky130_fd_sc_hd__a31o_2 _22892_ (.A1(_11471_),
    .A2(_12421_),
    .A3(_12423_),
    .B1(_05731_),
    .X(_12880_));
 sky130_fd_sc_hd__nor2_1 _22893_ (.A(net357),
    .B(_12880_),
    .Y(_12881_));
 sky130_fd_sc_hd__a21oi_2 _22894_ (.A1(_10963_),
    .A2(_10964_),
    .B1(_12880_),
    .Y(_12882_));
 sky130_fd_sc_hd__o21a_1 _22895_ (.A1(_10965_),
    .A2(_10967_),
    .B1(_12880_),
    .X(_12883_));
 sky130_fd_sc_hd__nor2_1 _22896_ (.A(_12882_),
    .B(_12883_),
    .Y(_12884_));
 sky130_fd_sc_hd__o21ai_1 _22897_ (.A1(_12433_),
    .A2(_12434_),
    .B1(_12430_),
    .Y(_12885_));
 sky130_fd_sc_hd__a21boi_2 _22898_ (.A1(_12430_),
    .A2(_12436_),
    .B1_N(_12884_),
    .Y(_12886_));
 sky130_fd_sc_hd__nand2_1 _22899_ (.A(_12885_),
    .B(_12884_),
    .Y(_12887_));
 sky130_fd_sc_hd__o221ai_4 _22900_ (.A1(_12882_),
    .A2(_12883_),
    .B1(_12433_),
    .B2(_12434_),
    .C1(_12430_),
    .Y(_12889_));
 sky130_fd_sc_hd__o21ai_1 _22901_ (.A1(_06793_),
    .A2(_06815_),
    .B1(_12889_),
    .Y(_12890_));
 sky130_fd_sc_hd__and3_1 _22902_ (.A(_06804_),
    .B(_06826_),
    .C(_12880_),
    .X(_12891_));
 sky130_fd_sc_hd__a21oi_1 _22903_ (.A1(_12887_),
    .A2(_12889_),
    .B1(_06848_),
    .Y(_12892_));
 sky130_fd_sc_hd__o22ai_4 _22904_ (.A1(net357),
    .A2(_12880_),
    .B1(_12886_),
    .B2(_12890_),
    .Y(_12893_));
 sky130_fd_sc_hd__inv_2 _22905_ (.A(_12893_),
    .Y(_12894_));
 sky130_fd_sc_hd__nor2_1 _22906_ (.A(net354),
    .B(_12894_),
    .Y(_12895_));
 sky130_fd_sc_hd__o21ai_4 _22907_ (.A1(_10487_),
    .A2(_10488_),
    .B1(_12893_),
    .Y(_12896_));
 sky130_fd_sc_hd__a31o_1 _22908_ (.A1(_12887_),
    .A2(_12889_),
    .A3(net357),
    .B1(_10492_),
    .X(_12897_));
 sky130_fd_sc_hd__o21ai_4 _22909_ (.A1(_12881_),
    .A2(_12897_),
    .B1(_12896_),
    .Y(_12898_));
 sky130_fd_sc_hd__a2bb2oi_4 _22910_ (.A1_N(_10026_),
    .A2_N(_12438_),
    .B1(_12445_),
    .B2(_12455_),
    .Y(_12900_));
 sky130_fd_sc_hd__o22ai_1 _22911_ (.A1(_10026_),
    .A2(_12438_),
    .B1(_12446_),
    .B2(_12456_),
    .Y(_12901_));
 sky130_fd_sc_hd__o211ai_2 _22912_ (.A1(_12897_),
    .A2(_12881_),
    .B1(_12896_),
    .C1(_12901_),
    .Y(_12902_));
 sky130_fd_sc_hd__o221a_1 _22913_ (.A1(_10026_),
    .A2(_12438_),
    .B1(_12446_),
    .B2(_12456_),
    .C1(_12898_),
    .X(_12903_));
 sky130_fd_sc_hd__o221ai_4 _22914_ (.A1(_10026_),
    .A2(_12438_),
    .B1(_12446_),
    .B2(_12456_),
    .C1(_12898_),
    .Y(_12904_));
 sky130_fd_sc_hd__o22ai_4 _22915_ (.A1(net374),
    .A2(_07702_),
    .B1(_12898_),
    .B2(_12900_),
    .Y(_12905_));
 sky130_fd_sc_hd__o22a_2 _22916_ (.A1(net354),
    .A2(_12894_),
    .B1(_12903_),
    .B2(_12905_),
    .X(_12906_));
 sky130_fd_sc_hd__o22ai_4 _22917_ (.A1(net354),
    .A2(_12894_),
    .B1(_12903_),
    .B2(_12905_),
    .Y(_12907_));
 sky130_fd_sc_hd__or3_1 _22918_ (.A(_08678_),
    .B(_08700_),
    .C(_12906_),
    .X(_12908_));
 sky130_fd_sc_hd__o21a_1 _22919_ (.A1(net170),
    .A2(net169),
    .B1(_12907_),
    .X(_12909_));
 sky130_fd_sc_hd__o21ai_4 _22920_ (.A1(net170),
    .A2(net169),
    .B1(_12907_),
    .Y(_12911_));
 sky130_fd_sc_hd__a31o_1 _22921_ (.A1(_12902_),
    .A2(_12904_),
    .A3(net354),
    .B1(net151),
    .X(_12912_));
 sky130_fd_sc_hd__a311o_2 _22922_ (.A1(_12902_),
    .A2(_12904_),
    .A3(net354),
    .B1(net151),
    .C1(_12895_),
    .X(_12913_));
 sky130_fd_sc_hd__o21ai_1 _22923_ (.A1(_12895_),
    .A2(_12912_),
    .B1(_12911_),
    .Y(_12914_));
 sky130_fd_sc_hd__and3_1 _22924_ (.A(_11547_),
    .B(_11549_),
    .C(_11059_),
    .X(_12915_));
 sky130_fd_sc_hd__nand3_1 _22925_ (.A(_12474_),
    .B(_12915_),
    .C(_12028_),
    .Y(_12916_));
 sky130_fd_sc_hd__a31oi_1 _22926_ (.A1(_12474_),
    .A2(_12915_),
    .A3(_12028_),
    .B1(_12475_),
    .Y(_12917_));
 sky130_fd_sc_hd__o211ai_4 _22927_ (.A1(_12473_),
    .A2(_12471_),
    .B1(_12916_),
    .C1(_12476_),
    .Y(_12918_));
 sky130_fd_sc_hd__nand4_1 _22928_ (.A(_12915_),
    .B(_12027_),
    .C(_12024_),
    .D(_11072_),
    .Y(_12919_));
 sky130_fd_sc_hd__nor3_1 _22929_ (.A(_12473_),
    .B(_12919_),
    .C(_12475_),
    .Y(_12920_));
 sky130_fd_sc_hd__nand3b_4 _22930_ (.A_N(_12919_),
    .B(_12476_),
    .C(_12474_),
    .Y(_12922_));
 sky130_fd_sc_hd__a22oi_2 _22931_ (.A1(_12911_),
    .A2(_12913_),
    .B1(_12918_),
    .B2(_12922_),
    .Y(_12923_));
 sky130_fd_sc_hd__a22o_1 _22932_ (.A1(_12911_),
    .A2(_12913_),
    .B1(_12918_),
    .B2(_12922_),
    .X(_12924_));
 sky130_fd_sc_hd__a211oi_2 _22933_ (.A1(_12477_),
    .A2(_12917_),
    .B1(_12920_),
    .C1(_12914_),
    .Y(_12925_));
 sky130_fd_sc_hd__nand4_4 _22934_ (.A(_12911_),
    .B(_12913_),
    .C(_12918_),
    .D(_12922_),
    .Y(_12926_));
 sky130_fd_sc_hd__nand3_2 _22935_ (.A(_12924_),
    .B(_12926_),
    .C(net338),
    .Y(_12927_));
 sky130_fd_sc_hd__o221a_1 _22936_ (.A1(net354),
    .A2(_12894_),
    .B1(_12903_),
    .B2(_12905_),
    .C1(_08732_),
    .X(_12928_));
 sky130_fd_sc_hd__a311o_1 _22937_ (.A1(_12902_),
    .A2(_12904_),
    .A3(net354),
    .B1(net338),
    .C1(_12895_),
    .X(_12929_));
 sky130_fd_sc_hd__a21oi_1 _22938_ (.A1(_12924_),
    .A2(_12926_),
    .B1(_08732_),
    .Y(_12930_));
 sky130_fd_sc_hd__o22ai_4 _22939_ (.A1(_08678_),
    .A2(_08700_),
    .B1(_12923_),
    .B2(_12925_),
    .Y(_12931_));
 sky130_fd_sc_hd__o31a_2 _22940_ (.A1(_08678_),
    .A2(_08700_),
    .A3(_12906_),
    .B1(_12927_),
    .X(_12933_));
 sky130_fd_sc_hd__o221ai_4 _22941_ (.A1(net174),
    .A2(_12480_),
    .B1(_12043_),
    .B2(_12048_),
    .C1(_12042_),
    .Y(_12934_));
 sky130_fd_sc_hd__o32a_1 _22942_ (.A1(_09134_),
    .A2(net193),
    .A3(_12481_),
    .B1(_12486_),
    .B2(_12482_),
    .X(_12935_));
 sky130_fd_sc_hd__a21oi_1 _22943_ (.A1(_12485_),
    .A2(_12934_),
    .B1(_09595_),
    .Y(_12936_));
 sky130_fd_sc_hd__a31oi_2 _22944_ (.A1(_09595_),
    .A2(_12485_),
    .A3(_12934_),
    .B1(_09840_),
    .Y(_12937_));
 sky130_fd_sc_hd__a31o_1 _22945_ (.A1(_09595_),
    .A2(_12485_),
    .A3(_12934_),
    .B1(_09840_),
    .X(_12938_));
 sky130_fd_sc_hd__o2111ai_4 _22946_ (.A1(_09595_),
    .A2(_12935_),
    .B1(_12931_),
    .C1(_12929_),
    .D1(_12937_),
    .Y(_12939_));
 sky130_fd_sc_hd__o21ai_1 _22947_ (.A1(_12936_),
    .A2(_12938_),
    .B1(_12933_),
    .Y(_12940_));
 sky130_fd_sc_hd__or4_2 _22948_ (.A(net351),
    .B(_09807_),
    .C(_12928_),
    .D(_12930_),
    .X(_12941_));
 sky130_fd_sc_hd__a2bb2oi_1 _22949_ (.A1_N(_09588_),
    .A2_N(net187),
    .B1(_12908_),
    .B2(_12927_),
    .Y(_12942_));
 sky130_fd_sc_hd__o221ai_4 _22950_ (.A1(_09588_),
    .A2(net187),
    .B1(_12907_),
    .B2(net338),
    .C1(_12931_),
    .Y(_12944_));
 sky130_fd_sc_hd__o211a_1 _22951_ (.A1(net338),
    .A2(_12906_),
    .B1(net172),
    .C1(_12927_),
    .X(_12945_));
 sky130_fd_sc_hd__o211ai_2 _22952_ (.A1(net338),
    .A2(_12906_),
    .B1(net172),
    .C1(_12927_),
    .Y(_12946_));
 sky130_fd_sc_hd__o2bb2ai_1 _22953_ (.A1_N(_12485_),
    .A2_N(_12934_),
    .B1(_12942_),
    .B2(_12945_),
    .Y(_12947_));
 sky130_fd_sc_hd__nand3_1 _22954_ (.A(_12935_),
    .B(_12944_),
    .C(_12946_),
    .Y(_12948_));
 sky130_fd_sc_hd__nand3_4 _22955_ (.A(_12947_),
    .B(_12948_),
    .C(net335),
    .Y(_12949_));
 sky130_fd_sc_hd__o21ai_4 _22956_ (.A1(net335),
    .A2(_12933_),
    .B1(_12949_),
    .Y(_12950_));
 sky130_fd_sc_hd__o211ai_4 _22957_ (.A1(_09134_),
    .A2(net193),
    .B1(_12939_),
    .C1(_12940_),
    .Y(_12951_));
 sky130_fd_sc_hd__o311a_1 _22958_ (.A1(net335),
    .A2(_12928_),
    .A3(_12930_),
    .B1(net174),
    .C1(_12949_),
    .X(_12952_));
 sky130_fd_sc_hd__nand3_4 _22959_ (.A(_12949_),
    .B(net174),
    .C(_12941_),
    .Y(_12953_));
 sky130_fd_sc_hd__o21ai_2 _22960_ (.A1(net177),
    .A2(_12495_),
    .B1(_12502_),
    .Y(_12955_));
 sky130_fd_sc_hd__a22oi_2 _22961_ (.A1(_12951_),
    .A2(_12953_),
    .B1(_12955_),
    .B2(_12500_),
    .Y(_12956_));
 sky130_fd_sc_hd__a22o_1 _22962_ (.A1(_12951_),
    .A2(_12953_),
    .B1(_12955_),
    .B2(_12500_),
    .X(_12957_));
 sky130_fd_sc_hd__o2111a_1 _22963_ (.A1(_12493_),
    .A2(net175),
    .B1(_12953_),
    .C1(_12951_),
    .D1(_12955_),
    .X(_12958_));
 sky130_fd_sc_hd__o2111ai_4 _22964_ (.A1(_12493_),
    .A2(net175),
    .B1(_12953_),
    .C1(_12951_),
    .D1(_12955_),
    .Y(_12959_));
 sky130_fd_sc_hd__o22ai_2 _22965_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_12956_),
    .B2(_12958_),
    .Y(_12960_));
 sky130_fd_sc_hd__a21o_1 _22966_ (.A1(_12941_),
    .A2(_12949_),
    .B1(net332),
    .X(_12961_));
 sky130_fd_sc_hd__inv_2 _22967_ (.A(_12961_),
    .Y(_12962_));
 sky130_fd_sc_hd__nand3_1 _22968_ (.A(_12957_),
    .B(_12959_),
    .C(net332),
    .Y(_12963_));
 sky130_fd_sc_hd__a31o_1 _22969_ (.A1(_12957_),
    .A2(_12959_),
    .A3(net332),
    .B1(_12962_),
    .X(_12964_));
 sky130_fd_sc_hd__o31a_2 _22970_ (.A1(_11079_),
    .A2(_12956_),
    .A3(_12958_),
    .B1(_12961_),
    .X(_12966_));
 sky130_fd_sc_hd__a2bb2oi_1 _22971_ (.A1_N(_08724_),
    .A2_N(_08726_),
    .B1(_12961_),
    .B2(_12963_),
    .Y(_12967_));
 sky130_fd_sc_hd__o221ai_4 _22972_ (.A1(_08724_),
    .A2(_08726_),
    .B1(_12950_),
    .B2(net332),
    .C1(_12960_),
    .Y(_12968_));
 sky130_fd_sc_hd__a311oi_2 _22973_ (.A1(_12957_),
    .A2(_12959_),
    .A3(net332),
    .B1(net175),
    .C1(_12962_),
    .Y(_12969_));
 sky130_fd_sc_hd__a311o_2 _22974_ (.A1(_12957_),
    .A2(_12959_),
    .A3(net332),
    .B1(net175),
    .C1(_12962_),
    .X(_12970_));
 sky130_fd_sc_hd__o2bb2ai_1 _22975_ (.A1_N(_12523_),
    .A2_N(_12525_),
    .B1(net199),
    .B2(_12511_),
    .Y(_12971_));
 sky130_fd_sc_hd__o211ai_1 _22976_ (.A1(net198),
    .A2(_12510_),
    .B1(_12523_),
    .C1(_12525_),
    .Y(_12972_));
 sky130_fd_sc_hd__o221ai_4 _22977_ (.A1(_12511_),
    .A2(net199),
    .B1(_12969_),
    .B2(_12967_),
    .C1(_12529_),
    .Y(_12973_));
 sky130_fd_sc_hd__o2111ai_4 _22978_ (.A1(net198),
    .A2(_12510_),
    .B1(_12968_),
    .C1(_12970_),
    .D1(_12971_),
    .Y(_12974_));
 sky130_fd_sc_hd__nand3_4 _22979_ (.A(_12973_),
    .B(_12974_),
    .C(net311),
    .Y(_12975_));
 sky130_fd_sc_hd__or3_2 _22980_ (.A(net329),
    .B(net327),
    .C(_12966_),
    .X(_12977_));
 sky130_fd_sc_hd__o31a_4 _22981_ (.A1(net329),
    .A2(net327),
    .A3(_12966_),
    .B1(_12975_),
    .X(_12978_));
 sky130_fd_sc_hd__a21oi_4 _22982_ (.A1(_12975_),
    .A2(_12977_),
    .B1(net308),
    .Y(_12979_));
 sky130_fd_sc_hd__or3_2 _22983_ (.A(_00011_),
    .B(net323),
    .C(_12978_),
    .X(_12980_));
 sky130_fd_sc_hd__a21oi_2 _22984_ (.A1(_12975_),
    .A2(_12977_),
    .B1(net199),
    .Y(_12981_));
 sky130_fd_sc_hd__a22o_1 _22985_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_12975_),
    .B2(_12977_),
    .X(_12982_));
 sky130_fd_sc_hd__a31oi_4 _22986_ (.A1(_12973_),
    .A2(_12974_),
    .A3(net311),
    .B1(net198),
    .Y(_12983_));
 sky130_fd_sc_hd__o21ai_4 _22987_ (.A1(net311),
    .A2(_12966_),
    .B1(_12983_),
    .Y(_12984_));
 sky130_fd_sc_hd__a21oi_2 _22988_ (.A1(_12977_),
    .A2(_12983_),
    .B1(_12981_),
    .Y(_12985_));
 sky130_fd_sc_hd__o2111a_1 _22989_ (.A1(_11138_),
    .A2(_11132_),
    .B1(_11136_),
    .C1(_11628_),
    .D1(_11629_),
    .X(_12986_));
 sky130_fd_sc_hd__o211a_2 _22990_ (.A1(_12079_),
    .A2(_12100_),
    .B1(_12986_),
    .C1(_12098_),
    .X(_12988_));
 sky130_fd_sc_hd__nand2_1 _22991_ (.A(_12988_),
    .B(_12540_),
    .Y(_12989_));
 sky130_fd_sc_hd__a32oi_4 _22992_ (.A1(_07936_),
    .A2(_12533_),
    .A3(_12534_),
    .B1(_12988_),
    .B2(_12540_),
    .Y(_12990_));
 sky130_fd_sc_hd__o211ai_4 _22993_ (.A1(_12539_),
    .A2(_12543_),
    .B1(_12989_),
    .C1(_12537_),
    .Y(_12991_));
 sky130_fd_sc_hd__o211ai_4 _22994_ (.A1(_11147_),
    .A2(_11149_),
    .B1(_12988_),
    .C1(_12537_),
    .Y(_12992_));
 sky130_fd_sc_hd__nand4_1 _22995_ (.A(_12537_),
    .B(_12988_),
    .C(_12540_),
    .D(_11150_),
    .Y(_12993_));
 sky130_fd_sc_hd__a2bb2oi_4 _22996_ (.A1_N(_12539_),
    .A2_N(_12992_),
    .B1(_12545_),
    .B2(_12990_),
    .Y(_12994_));
 sky130_fd_sc_hd__o2111a_2 _22997_ (.A1(_12992_),
    .A2(_12539_),
    .B1(_12984_),
    .C1(_12991_),
    .D1(_12982_),
    .X(_12995_));
 sky130_fd_sc_hd__o2111ai_4 _22998_ (.A1(_12992_),
    .A2(_12539_),
    .B1(_12984_),
    .C1(_12991_),
    .D1(_12982_),
    .Y(_12996_));
 sky130_fd_sc_hd__a22o_2 _22999_ (.A1(_12982_),
    .A2(_12984_),
    .B1(_12991_),
    .B2(_12993_),
    .X(_12997_));
 sky130_fd_sc_hd__o22ai_4 _23000_ (.A1(_00011_),
    .A2(net321),
    .B1(_12985_),
    .B2(_12994_),
    .Y(_12999_));
 sky130_fd_sc_hd__o211ai_4 _23001_ (.A1(_00011_),
    .A2(net323),
    .B1(_12996_),
    .C1(_12997_),
    .Y(_13000_));
 sky130_fd_sc_hd__a31oi_4 _23002_ (.A1(_12997_),
    .A2(net307),
    .A3(_12996_),
    .B1(_12979_),
    .Y(_13001_));
 sky130_fd_sc_hd__o22ai_4 _23003_ (.A1(net307),
    .A2(_12978_),
    .B1(_12995_),
    .B2(_12999_),
    .Y(_13002_));
 sky130_fd_sc_hd__a21oi_4 _23004_ (.A1(_12980_),
    .A2(_13000_),
    .B1(net278),
    .Y(_13003_));
 sky130_fd_sc_hd__or3_2 _23005_ (.A(net304),
    .B(_01951_),
    .C(_13001_),
    .X(_13004_));
 sky130_fd_sc_hd__a311oi_4 _23006_ (.A1(_12997_),
    .A2(net307),
    .A3(_12996_),
    .B1(_07936_),
    .C1(_12979_),
    .Y(_13005_));
 sky130_fd_sc_hd__o221ai_4 _23007_ (.A1(net307),
    .A2(_12978_),
    .B1(_12995_),
    .B2(_12999_),
    .C1(_07935_),
    .Y(_13006_));
 sky130_fd_sc_hd__a2bb2oi_2 _23008_ (.A1_N(_07928_),
    .A2_N(_07930_),
    .B1(_12980_),
    .B2(_13000_),
    .Y(_13007_));
 sky130_fd_sc_hd__o21ai_4 _23009_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_13002_),
    .Y(_13008_));
 sky130_fd_sc_hd__o32a_1 _23010_ (.A1(_07555_),
    .A2(_07557_),
    .A3(_12547_),
    .B1(_12552_),
    .B2(_12548_),
    .X(_13010_));
 sky130_fd_sc_hd__o32ai_4 _23011_ (.A1(_07555_),
    .A2(_07557_),
    .A3(_12547_),
    .B1(_12552_),
    .B2(_12548_),
    .Y(_13011_));
 sky130_fd_sc_hd__o21ai_4 _23012_ (.A1(_13005_),
    .A2(_13007_),
    .B1(_13011_),
    .Y(_13012_));
 sky130_fd_sc_hd__nand3_4 _23013_ (.A(_13010_),
    .B(_13008_),
    .C(_13006_),
    .Y(_13013_));
 sky130_fd_sc_hd__o311a_1 _23014_ (.A1(_13005_),
    .A2(_13007_),
    .A3(_13011_),
    .B1(net278),
    .C1(_13012_),
    .X(_13014_));
 sky130_fd_sc_hd__nand3_2 _23015_ (.A(_13012_),
    .B(_13013_),
    .C(net279),
    .Y(_13015_));
 sky130_fd_sc_hd__a31o_2 _23016_ (.A1(_13012_),
    .A2(_13013_),
    .A3(net278),
    .B1(_13003_),
    .X(_13016_));
 sky130_fd_sc_hd__o221a_1 _23017_ (.A1(net227),
    .A2(_12120_),
    .B1(_12559_),
    .B2(net224),
    .C1(_12565_),
    .X(_13017_));
 sky130_fd_sc_hd__o221ai_4 _23018_ (.A1(net227),
    .A2(_12120_),
    .B1(_12559_),
    .B2(net224),
    .C1(_12565_),
    .Y(_13018_));
 sky130_fd_sc_hd__a22oi_2 _23019_ (.A1(net224),
    .A2(_12559_),
    .B1(_12565_),
    .B2(_12125_),
    .Y(_13019_));
 sky130_fd_sc_hd__a31oi_2 _23020_ (.A1(_13012_),
    .A2(_13013_),
    .A3(net278),
    .B1(net202),
    .Y(_13021_));
 sky130_fd_sc_hd__a311oi_4 _23021_ (.A1(_13012_),
    .A2(_13013_),
    .A3(net278),
    .B1(net202),
    .C1(_13003_),
    .Y(_13022_));
 sky130_fd_sc_hd__o211ai_4 _23022_ (.A1(net279),
    .A2(_13001_),
    .B1(_07564_),
    .C1(_13015_),
    .Y(_13023_));
 sky130_fd_sc_hd__a2bb2oi_4 _23023_ (.A1_N(_07555_),
    .A2_N(_07557_),
    .B1(_13004_),
    .B2(_13015_),
    .Y(_13024_));
 sky130_fd_sc_hd__o22ai_2 _23024_ (.A1(_07555_),
    .A2(_07557_),
    .B1(_13003_),
    .B2(_13014_),
    .Y(_13025_));
 sky130_fd_sc_hd__a21oi_1 _23025_ (.A1(_13004_),
    .A2(_13021_),
    .B1(_13024_),
    .Y(_13026_));
 sky130_fd_sc_hd__o211ai_2 _23026_ (.A1(_12563_),
    .A2(_13017_),
    .B1(_13023_),
    .C1(_13025_),
    .Y(_13027_));
 sky130_fd_sc_hd__o22ai_2 _23027_ (.A1(_12561_),
    .A2(_13019_),
    .B1(_13022_),
    .B2(_13024_),
    .Y(_13028_));
 sky130_fd_sc_hd__nand3_4 _23028_ (.A(_13027_),
    .B(_13028_),
    .C(net277),
    .Y(_13029_));
 sky130_fd_sc_hd__o22a_1 _23029_ (.A1(_03986_),
    .A2(_03997_),
    .B1(_13003_),
    .B2(_13014_),
    .X(_13030_));
 sky130_fd_sc_hd__inv_2 _23030_ (.A(_13030_),
    .Y(_13032_));
 sky130_fd_sc_hd__o211ai_1 _23031_ (.A1(_12561_),
    .A2(_13019_),
    .B1(_13023_),
    .C1(_13025_),
    .Y(_13033_));
 sky130_fd_sc_hd__o22ai_1 _23032_ (.A1(_12563_),
    .A2(_13017_),
    .B1(_13022_),
    .B2(_13024_),
    .Y(_13034_));
 sky130_fd_sc_hd__nand3_1 _23033_ (.A(_13033_),
    .B(_13034_),
    .C(net277),
    .Y(_13035_));
 sky130_fd_sc_hd__o21ai_4 _23034_ (.A1(net277),
    .A2(_13016_),
    .B1(_13029_),
    .Y(_13036_));
 sky130_fd_sc_hd__o311a_1 _23035_ (.A1(net277),
    .A2(_13003_),
    .A3(_13014_),
    .B1(_13029_),
    .C1(net222),
    .X(_13037_));
 sky130_fd_sc_hd__o211ai_4 _23036_ (.A1(_13016_),
    .A2(net277),
    .B1(net222),
    .C1(_13029_),
    .Y(_13038_));
 sky130_fd_sc_hd__nand3_4 _23037_ (.A(_13035_),
    .B(net224),
    .C(_13032_),
    .Y(_13039_));
 sky130_fd_sc_hd__nand2_1 _23038_ (.A(_13038_),
    .B(_13039_),
    .Y(_13040_));
 sky130_fd_sc_hd__a22o_1 _23039_ (.A1(net225),
    .A2(_12573_),
    .B1(_12587_),
    .B2(_12590_),
    .X(_13041_));
 sky130_fd_sc_hd__o211ai_4 _23040_ (.A1(_12578_),
    .A2(_12570_),
    .B1(_12590_),
    .C1(_12587_),
    .Y(_13043_));
 sky130_fd_sc_hd__a31oi_2 _23041_ (.A1(_12580_),
    .A2(_12587_),
    .A3(_12590_),
    .B1(_12575_),
    .Y(_13044_));
 sky130_fd_sc_hd__o2111ai_4 _23042_ (.A1(net225),
    .A2(_12573_),
    .B1(_13038_),
    .C1(_13039_),
    .D1(_13041_),
    .Y(_13045_));
 sky130_fd_sc_hd__a22oi_4 _23043_ (.A1(_13038_),
    .A2(_13039_),
    .B1(_13041_),
    .B2(_12580_),
    .Y(_13046_));
 sky130_fd_sc_hd__o211ai_2 _23044_ (.A1(net227),
    .A2(_12572_),
    .B1(_12596_),
    .C1(_13040_),
    .Y(_13047_));
 sky130_fd_sc_hd__o21ai_4 _23045_ (.A1(_13040_),
    .A2(_13044_),
    .B1(net272),
    .Y(_13048_));
 sky130_fd_sc_hd__nand3_1 _23046_ (.A(_13045_),
    .B(_13047_),
    .C(net272),
    .Y(_13049_));
 sky130_fd_sc_hd__o311a_1 _23047_ (.A1(net277),
    .A2(_13003_),
    .A3(_13014_),
    .B1(_13029_),
    .C1(_05234_),
    .X(_13050_));
 sky130_fd_sc_hd__or3_2 _23048_ (.A(net296),
    .B(_05232_),
    .C(_13036_),
    .X(_13051_));
 sky130_fd_sc_hd__o32a_2 _23049_ (.A1(net296),
    .A2(_05232_),
    .A3(_13036_),
    .B1(_13046_),
    .B2(_13048_),
    .X(_13052_));
 sky130_fd_sc_hd__o22ai_4 _23050_ (.A1(net272),
    .A2(_13036_),
    .B1(_13046_),
    .B2(_13048_),
    .Y(_13054_));
 sky130_fd_sc_hd__a22oi_4 _23051_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_13049_),
    .B2(_13051_),
    .Y(_13055_));
 sky130_fd_sc_hd__o21ai_4 _23052_ (.A1(_06914_),
    .A2(net250),
    .B1(_13054_),
    .Y(_13056_));
 sky130_fd_sc_hd__a31oi_1 _23053_ (.A1(_13045_),
    .A2(_13047_),
    .A3(net272),
    .B1(net225),
    .Y(_13057_));
 sky130_fd_sc_hd__a311oi_2 _23054_ (.A1(_13045_),
    .A2(_13047_),
    .A3(net272),
    .B1(_13050_),
    .C1(net225),
    .Y(_13058_));
 sky130_fd_sc_hd__o221ai_4 _23055_ (.A1(net272),
    .A2(_13036_),
    .B1(_13046_),
    .B2(_13048_),
    .C1(net227),
    .Y(_13059_));
 sky130_fd_sc_hd__a21oi_2 _23056_ (.A1(_13051_),
    .A2(_13057_),
    .B1(_13055_),
    .Y(_13060_));
 sky130_fd_sc_hd__nand2_1 _23057_ (.A(_13056_),
    .B(_13059_),
    .Y(_13061_));
 sky130_fd_sc_hd__and4_1 _23058_ (.A(_11212_),
    .B(_11213_),
    .C(_11701_),
    .D(_11703_),
    .X(_13062_));
 sky130_fd_sc_hd__nand4_1 _23059_ (.A(_11212_),
    .B(_11213_),
    .C(_11701_),
    .D(_11703_),
    .Y(_13063_));
 sky130_fd_sc_hd__a211oi_2 _23060_ (.A1(_12149_),
    .A2(_12169_),
    .B1(_13063_),
    .C1(_12172_),
    .Y(_13065_));
 sky130_fd_sc_hd__nand3_2 _23061_ (.A(_12606_),
    .B(_13062_),
    .C(_12174_),
    .Y(_13066_));
 sky130_fd_sc_hd__a32oi_1 _23062_ (.A1(net232),
    .A2(_12574_),
    .A3(_12598_),
    .B1(_13065_),
    .B2(_12606_),
    .Y(_13067_));
 sky130_fd_sc_hd__o211a_2 _23063_ (.A1(_12610_),
    .A2(_12605_),
    .B1(_12607_),
    .C1(_13066_),
    .X(_13068_));
 sky130_fd_sc_hd__o211ai_4 _23064_ (.A1(_12610_),
    .A2(_12605_),
    .B1(_12607_),
    .C1(_13066_),
    .Y(_13069_));
 sky130_fd_sc_hd__nand4_1 _23065_ (.A(_12606_),
    .B(_12607_),
    .C(_13062_),
    .D(_12174_),
    .Y(_13070_));
 sky130_fd_sc_hd__nand4_1 _23066_ (.A(_12607_),
    .B(_13062_),
    .C(_11224_),
    .D(_12174_),
    .Y(_13071_));
 sky130_fd_sc_hd__nand4_4 _23067_ (.A(_12606_),
    .B(_13065_),
    .C(_12607_),
    .D(_11224_),
    .Y(_13072_));
 sky130_fd_sc_hd__inv_2 _23068_ (.A(_13072_),
    .Y(_13073_));
 sky130_fd_sc_hd__a2bb2oi_1 _23069_ (.A1_N(_12605_),
    .A2_N(_13071_),
    .B1(_12612_),
    .B2(_13067_),
    .Y(_13074_));
 sky130_fd_sc_hd__a31o_1 _23070_ (.A1(_12607_),
    .A2(_12612_),
    .A3(_13066_),
    .B1(_13073_),
    .X(_13076_));
 sky130_fd_sc_hd__a21oi_2 _23071_ (.A1(_13069_),
    .A2(_13072_),
    .B1(_13061_),
    .Y(_13077_));
 sky130_fd_sc_hd__o221ai_2 _23072_ (.A1(_11225_),
    .A2(_13070_),
    .B1(_13058_),
    .B2(_13055_),
    .C1(_13069_),
    .Y(_13078_));
 sky130_fd_sc_hd__o21ai_2 _23073_ (.A1(net270),
    .A2(_05483_),
    .B1(_13078_),
    .Y(_13079_));
 sky130_fd_sc_hd__nand4_4 _23074_ (.A(_13056_),
    .B(_13059_),
    .C(_13069_),
    .D(_13072_),
    .Y(_13080_));
 sky130_fd_sc_hd__a22o_1 _23075_ (.A1(_13056_),
    .A2(_13059_),
    .B1(_13069_),
    .B2(_13072_),
    .X(_13081_));
 sky130_fd_sc_hd__o221ai_4 _23076_ (.A1(net270),
    .A2(_05483_),
    .B1(_13060_),
    .B2(_13074_),
    .C1(_13080_),
    .Y(_13082_));
 sky130_fd_sc_hd__a211o_1 _23077_ (.A1(_13049_),
    .A2(_13051_),
    .B1(net270),
    .C1(net268),
    .X(_13083_));
 sky130_fd_sc_hd__inv_2 _23078_ (.A(_13083_),
    .Y(_13084_));
 sky130_fd_sc_hd__a31o_1 _23079_ (.A1(_13081_),
    .A2(net245),
    .A3(_13080_),
    .B1(_13084_),
    .X(_13085_));
 sky130_fd_sc_hd__a311oi_4 _23080_ (.A1(_13081_),
    .A2(net245),
    .A3(_13080_),
    .B1(_13084_),
    .C1(net232),
    .Y(_13087_));
 sky130_fd_sc_hd__o211ai_4 _23081_ (.A1(net245),
    .A2(_13052_),
    .B1(net234),
    .C1(_13082_),
    .Y(_13088_));
 sky130_fd_sc_hd__a21oi_1 _23082_ (.A1(_13082_),
    .A2(_13083_),
    .B1(net234),
    .Y(_13089_));
 sky130_fd_sc_hd__o221ai_4 _23083_ (.A1(net245),
    .A2(_13054_),
    .B1(_13077_),
    .B2(_13079_),
    .C1(net233),
    .Y(_13090_));
 sky130_fd_sc_hd__o221a_1 _23084_ (.A1(_12190_),
    .A2(_12185_),
    .B1(_06314_),
    .B2(_12614_),
    .C1(_12183_),
    .X(_13091_));
 sky130_fd_sc_hd__o21ai_1 _23085_ (.A1(_06314_),
    .A2(_12614_),
    .B1(_12619_),
    .Y(_13092_));
 sky130_fd_sc_hd__o21ai_2 _23086_ (.A1(_12621_),
    .A2(_12619_),
    .B1(_12624_),
    .Y(_13093_));
 sky130_fd_sc_hd__a21oi_2 _23087_ (.A1(_12622_),
    .A2(_12618_),
    .B1(_12623_),
    .Y(_13094_));
 sky130_fd_sc_hd__a21oi_1 _23088_ (.A1(_13088_),
    .A2(_13090_),
    .B1(_13093_),
    .Y(_13095_));
 sky130_fd_sc_hd__o2bb2ai_4 _23089_ (.A1_N(_13088_),
    .A2_N(_13090_),
    .B1(_13091_),
    .B2(_12621_),
    .Y(_13096_));
 sky130_fd_sc_hd__o2111a_1 _23090_ (.A1(net252),
    .A2(_12616_),
    .B1(_13088_),
    .C1(_13090_),
    .D1(_13092_),
    .X(_13098_));
 sky130_fd_sc_hd__nand3_4 _23091_ (.A(_13088_),
    .B(_13090_),
    .C(_13093_),
    .Y(_13099_));
 sky130_fd_sc_hd__o311a_1 _23092_ (.A1(_13094_),
    .A2(_13089_),
    .A3(_13087_),
    .B1(net242),
    .C1(_13096_),
    .X(_13100_));
 sky130_fd_sc_hd__nand3_1 _23093_ (.A(_13096_),
    .B(_13099_),
    .C(net242),
    .Y(_13101_));
 sky130_fd_sc_hd__o221a_4 _23094_ (.A1(net245),
    .A2(_13054_),
    .B1(_13077_),
    .B2(_13079_),
    .C1(_05754_),
    .X(_13102_));
 sky130_fd_sc_hd__a211o_1 _23095_ (.A1(_13082_),
    .A2(_13083_),
    .B1(_05750_),
    .C1(net264),
    .X(_13103_));
 sky130_fd_sc_hd__o22ai_2 _23096_ (.A1(_05750_),
    .A2(net264),
    .B1(_13095_),
    .B2(_13098_),
    .Y(_13104_));
 sky130_fd_sc_hd__a31oi_2 _23097_ (.A1(_13096_),
    .A2(_13099_),
    .A3(net242),
    .B1(_13102_),
    .Y(_13105_));
 sky130_fd_sc_hd__a31o_1 _23098_ (.A1(_13096_),
    .A2(_13099_),
    .A3(net242),
    .B1(net252),
    .X(_13106_));
 sky130_fd_sc_hd__a311oi_4 _23099_ (.A1(_13096_),
    .A2(_13099_),
    .A3(net242),
    .B1(_13102_),
    .C1(net252),
    .Y(_13107_));
 sky130_fd_sc_hd__a311o_1 _23100_ (.A1(_13096_),
    .A2(_13099_),
    .A3(net242),
    .B1(_13102_),
    .C1(net252),
    .X(_13109_));
 sky130_fd_sc_hd__a21oi_4 _23101_ (.A1(_13101_),
    .A2(_13103_),
    .B1(_06314_),
    .Y(_13110_));
 sky130_fd_sc_hd__o221ai_4 _23102_ (.A1(net284),
    .A2(_06307_),
    .B1(_13085_),
    .B2(net242),
    .C1(_13104_),
    .Y(_13111_));
 sky130_fd_sc_hd__a31oi_4 _23103_ (.A1(_12201_),
    .A2(_12219_),
    .A3(_12635_),
    .B1(_12636_),
    .Y(_13112_));
 sky130_fd_sc_hd__a31o_1 _23104_ (.A1(_12201_),
    .A2(_12219_),
    .A3(_12635_),
    .B1(_12636_),
    .X(_13113_));
 sky130_fd_sc_hd__nand3_1 _23105_ (.A(_13109_),
    .B(_13111_),
    .C(_13113_),
    .Y(_13114_));
 sky130_fd_sc_hd__o21ai_1 _23106_ (.A1(_13107_),
    .A2(_13110_),
    .B1(_13112_),
    .Y(_13115_));
 sky130_fd_sc_hd__o211ai_2 _23107_ (.A1(net260),
    .A2(net258),
    .B1(_13114_),
    .C1(_13115_),
    .Y(_13116_));
 sky130_fd_sc_hd__o311a_2 _23108_ (.A1(_05750_),
    .A2(net264),
    .A3(_13085_),
    .B1(_05995_),
    .C1(_13104_),
    .X(_13117_));
 sky130_fd_sc_hd__or3_1 _23109_ (.A(net260),
    .B(net258),
    .C(_13105_),
    .X(_13118_));
 sky130_fd_sc_hd__o21ai_2 _23110_ (.A1(_13107_),
    .A2(_13110_),
    .B1(_13113_),
    .Y(_13120_));
 sky130_fd_sc_hd__o21ai_1 _23111_ (.A1(_06314_),
    .A2(_13105_),
    .B1(_13112_),
    .Y(_13121_));
 sky130_fd_sc_hd__o211ai_4 _23112_ (.A1(_13102_),
    .A2(_13106_),
    .B1(_13112_),
    .C1(_13111_),
    .Y(_13122_));
 sky130_fd_sc_hd__o221ai_2 _23113_ (.A1(net260),
    .A2(net258),
    .B1(_13107_),
    .B2(_13121_),
    .C1(_13120_),
    .Y(_13123_));
 sky130_fd_sc_hd__a31oi_4 _23114_ (.A1(net240),
    .A2(_13120_),
    .A3(_13122_),
    .B1(_13117_),
    .Y(_13124_));
 sky130_fd_sc_hd__a311o_1 _23115_ (.A1(net240),
    .A2(_13120_),
    .A3(_13122_),
    .B1(net213),
    .C1(_13117_),
    .X(_13125_));
 sky130_fd_sc_hd__a2bb2oi_1 _23116_ (.A1_N(_06009_),
    .A2_N(net287),
    .B1(_13118_),
    .B2(_13123_),
    .Y(_13126_));
 sky130_fd_sc_hd__o311ai_4 _23117_ (.A1(net240),
    .A2(_13100_),
    .A3(_13102_),
    .B1(_13116_),
    .C1(_06014_),
    .Y(_13127_));
 sky130_fd_sc_hd__o221a_2 _23118_ (.A1(_06011_),
    .A2(_06012_),
    .B1(_13105_),
    .B2(net240),
    .C1(_13123_),
    .X(_13128_));
 sky130_fd_sc_hd__a311o_1 _23119_ (.A1(net240),
    .A2(_13120_),
    .A3(_13122_),
    .B1(_06014_),
    .C1(_13117_),
    .X(_13129_));
 sky130_fd_sc_hd__a31o_1 _23120_ (.A1(_12655_),
    .A2(_12661_),
    .A3(_12663_),
    .B1(_12652_),
    .X(_13131_));
 sky130_fd_sc_hd__a31oi_1 _23121_ (.A1(_12655_),
    .A2(_12661_),
    .A3(_12663_),
    .B1(_12652_),
    .Y(_13132_));
 sky130_fd_sc_hd__o2111ai_1 _23122_ (.A1(net263),
    .A2(_12650_),
    .B1(_12671_),
    .C1(_13127_),
    .D1(_13129_),
    .Y(_13133_));
 sky130_fd_sc_hd__o21ai_1 _23123_ (.A1(_13126_),
    .A2(_13128_),
    .B1(_13131_),
    .Y(_13134_));
 sky130_fd_sc_hd__nand3_1 _23124_ (.A(_13134_),
    .B(net213),
    .C(_13133_),
    .Y(_13135_));
 sky130_fd_sc_hd__or3_1 _23125_ (.A(net239),
    .B(_06292_),
    .C(_13124_),
    .X(_13136_));
 sky130_fd_sc_hd__o21ai_1 _23126_ (.A1(_13126_),
    .A2(_13128_),
    .B1(_13132_),
    .Y(_13137_));
 sky130_fd_sc_hd__nand3_2 _23127_ (.A(_13131_),
    .B(_13129_),
    .C(_13127_),
    .Y(_13138_));
 sky130_fd_sc_hd__o211ai_4 _23128_ (.A1(net239),
    .A2(_06292_),
    .B1(_13137_),
    .C1(_13138_),
    .Y(_13139_));
 sky130_fd_sc_hd__o21ai_4 _23129_ (.A1(net213),
    .A2(_13124_),
    .B1(_13139_),
    .Y(_13140_));
 sky130_fd_sc_hd__o31a_2 _23130_ (.A1(net239),
    .A2(_06292_),
    .A3(_13124_),
    .B1(_13139_),
    .X(_13142_));
 sky130_fd_sc_hd__nand3_4 _23131_ (.A(net261),
    .B(_13125_),
    .C(_13135_),
    .Y(_13143_));
 sky130_fd_sc_hd__nand3_1 _23132_ (.A(_13139_),
    .B(net263),
    .C(_13136_),
    .Y(_13144_));
 sky130_fd_sc_hd__nand2_1 _23133_ (.A(_13143_),
    .B(_13144_),
    .Y(_13145_));
 sky130_fd_sc_hd__and4_1 _23134_ (.A(_11289_),
    .B(_11291_),
    .C(_11778_),
    .D(_11780_),
    .X(_13146_));
 sky130_fd_sc_hd__nor3b_1 _23135_ (.A(_12244_),
    .B(_12246_),
    .C_N(_13146_),
    .Y(_13147_));
 sky130_fd_sc_hd__nand3_1 _23136_ (.A(_12675_),
    .B(_13146_),
    .C(_12248_),
    .Y(_13148_));
 sky130_fd_sc_hd__o211ai_4 _23137_ (.A1(_12679_),
    .A2(_12674_),
    .B1(_12676_),
    .C1(_13148_),
    .Y(_13149_));
 sky130_fd_sc_hd__nand4_4 _23138_ (.A(_12675_),
    .B(_13147_),
    .C(_12676_),
    .D(_11300_),
    .Y(_13150_));
 sky130_fd_sc_hd__nand2_1 _23139_ (.A(_13149_),
    .B(_13150_),
    .Y(_13151_));
 sky130_fd_sc_hd__a21oi_2 _23140_ (.A1(_13149_),
    .A2(_13150_),
    .B1(_13145_),
    .Y(_13153_));
 sky130_fd_sc_hd__a31o_1 _23141_ (.A1(_13145_),
    .A2(_13149_),
    .A3(_13150_),
    .B1(_06613_),
    .X(_13154_));
 sky130_fd_sc_hd__and3_1 _23142_ (.A(_06613_),
    .B(_13125_),
    .C(_13135_),
    .X(_13155_));
 sky130_fd_sc_hd__or3_2 _23143_ (.A(net238),
    .B(_06610_),
    .C(_13142_),
    .X(_13156_));
 sky130_fd_sc_hd__a22o_1 _23144_ (.A1(_13143_),
    .A2(_13144_),
    .B1(_13149_),
    .B2(_13150_),
    .X(_13157_));
 sky130_fd_sc_hd__o211ai_4 _23145_ (.A1(_13140_),
    .A2(net261),
    .B1(_13150_),
    .C1(_13149_),
    .Y(_13158_));
 sky130_fd_sc_hd__o2111ai_4 _23146_ (.A1(_05768_),
    .A2(_13140_),
    .B1(_13143_),
    .C1(_13149_),
    .D1(_13150_),
    .Y(_13159_));
 sky130_fd_sc_hd__nand3_2 _23147_ (.A(_13157_),
    .B(_13159_),
    .C(net210),
    .Y(_13160_));
 sky130_fd_sc_hd__o221a_4 _23148_ (.A1(net210),
    .A2(_13140_),
    .B1(_13153_),
    .B2(_13154_),
    .C1(_06904_),
    .X(_13161_));
 sky130_fd_sc_hd__a211o_1 _23149_ (.A1(_13156_),
    .A2(_13160_),
    .B1(_06899_),
    .C1(net228),
    .X(_13162_));
 sky130_fd_sc_hd__a311oi_4 _23150_ (.A1(_13157_),
    .A2(_13159_),
    .A3(net210),
    .B1(_13155_),
    .C1(net292),
    .Y(_13164_));
 sky130_fd_sc_hd__nand3_4 _23151_ (.A(_13160_),
    .B(_05507_),
    .C(_13156_),
    .Y(_13165_));
 sky130_fd_sc_hd__o221ai_4 _23152_ (.A1(net210),
    .A2(_13140_),
    .B1(_13153_),
    .B2(_13154_),
    .C1(net292),
    .Y(_13166_));
 sky130_fd_sc_hd__o221a_1 _23153_ (.A1(_12257_),
    .A2(net299),
    .B1(net295),
    .B2(_12686_),
    .C1(_12690_),
    .X(_13167_));
 sky130_fd_sc_hd__o221ai_4 _23154_ (.A1(_12257_),
    .A2(net299),
    .B1(net295),
    .B2(_12686_),
    .C1(_12690_),
    .Y(_13168_));
 sky130_fd_sc_hd__o22a_1 _23155_ (.A1(_12693_),
    .A2(_12684_),
    .B1(_12691_),
    .B2(_12695_),
    .X(_13169_));
 sky130_fd_sc_hd__o21ai_2 _23156_ (.A1(_12684_),
    .A2(_12693_),
    .B1(_13168_),
    .Y(_13170_));
 sky130_fd_sc_hd__a21oi_1 _23157_ (.A1(_13165_),
    .A2(_13166_),
    .B1(_13169_),
    .Y(_13171_));
 sky130_fd_sc_hd__o2bb2ai_4 _23158_ (.A1_N(_13165_),
    .A2_N(_13166_),
    .B1(_13167_),
    .B2(_12694_),
    .Y(_13172_));
 sky130_fd_sc_hd__o2111a_1 _23159_ (.A1(net294),
    .A2(_12687_),
    .B1(_13165_),
    .C1(_13166_),
    .D1(_13168_),
    .X(_13173_));
 sky130_fd_sc_hd__nand3_4 _23160_ (.A(_13165_),
    .B(_13166_),
    .C(_13169_),
    .Y(_13175_));
 sky130_fd_sc_hd__nand3_1 _23161_ (.A(_13172_),
    .B(_13175_),
    .C(net208),
    .Y(_13176_));
 sky130_fd_sc_hd__a311o_1 _23162_ (.A1(_13157_),
    .A2(_13159_),
    .A3(net210),
    .B1(net208),
    .C1(_13155_),
    .X(_13177_));
 sky130_fd_sc_hd__o22ai_2 _23163_ (.A1(_06899_),
    .A2(_06901_),
    .B1(_13171_),
    .B2(_13173_),
    .Y(_13178_));
 sky130_fd_sc_hd__a31oi_4 _23164_ (.A1(_13172_),
    .A2(_13175_),
    .A3(net208),
    .B1(_13161_),
    .Y(_13179_));
 sky130_fd_sc_hd__a31o_1 _23165_ (.A1(_13172_),
    .A2(_13175_),
    .A3(net208),
    .B1(_13161_),
    .X(_13180_));
 sky130_fd_sc_hd__a311o_1 _23166_ (.A1(_13172_),
    .A2(_13175_),
    .A3(net208),
    .B1(net185),
    .C1(_13161_),
    .X(_13181_));
 sky130_fd_sc_hd__o311a_1 _23167_ (.A1(_02093_),
    .A2(_02115_),
    .A3(_12271_),
    .B1(_12280_),
    .C1(_12707_),
    .X(_13182_));
 sky130_fd_sc_hd__o21ai_2 _23168_ (.A1(_12708_),
    .A2(_12712_),
    .B1(_12707_),
    .Y(_13183_));
 sky130_fd_sc_hd__a31oi_1 _23169_ (.A1(_13172_),
    .A2(_13175_),
    .A3(net208),
    .B1(net294),
    .Y(_13184_));
 sky130_fd_sc_hd__a311oi_4 _23170_ (.A1(_13172_),
    .A2(_13175_),
    .A3(net208),
    .B1(_13161_),
    .C1(net294),
    .Y(_13186_));
 sky130_fd_sc_hd__a311o_1 _23171_ (.A1(_13172_),
    .A2(_13175_),
    .A3(net208),
    .B1(_13161_),
    .C1(net294),
    .X(_13187_));
 sky130_fd_sc_hd__a2bb2oi_2 _23172_ (.A1_N(net318),
    .A2_N(net316),
    .B1(_13162_),
    .B2(_13176_),
    .Y(_13188_));
 sky130_fd_sc_hd__o211ai_2 _23173_ (.A1(net318),
    .A2(net316),
    .B1(_13177_),
    .C1(_13178_),
    .Y(_13189_));
 sky130_fd_sc_hd__o211ai_1 _23174_ (.A1(_12708_),
    .A2(_13182_),
    .B1(_13187_),
    .C1(_13189_),
    .Y(_13190_));
 sky130_fd_sc_hd__o21ai_1 _23175_ (.A1(_13186_),
    .A2(_13188_),
    .B1(_13183_),
    .Y(_13191_));
 sky130_fd_sc_hd__o211ai_2 _23176_ (.A1(_07227_),
    .A2(net206),
    .B1(_13190_),
    .C1(_13191_),
    .Y(_13192_));
 sky130_fd_sc_hd__or3_1 _23177_ (.A(_07227_),
    .B(_07229_),
    .C(_13179_),
    .X(_13193_));
 sky130_fd_sc_hd__o21ai_1 _23178_ (.A1(net295),
    .A2(_13179_),
    .B1(_13183_),
    .Y(_13194_));
 sky130_fd_sc_hd__o22ai_2 _23179_ (.A1(_12708_),
    .A2(_13182_),
    .B1(_13186_),
    .B2(_13188_),
    .Y(_13195_));
 sky130_fd_sc_hd__o221ai_4 _23180_ (.A1(_07227_),
    .A2(net206),
    .B1(_13186_),
    .B2(_13194_),
    .C1(_13195_),
    .Y(_13197_));
 sky130_fd_sc_hd__o21ai_2 _23181_ (.A1(net185),
    .A2(_13179_),
    .B1(_13197_),
    .Y(_13198_));
 sky130_fd_sc_hd__or3_2 _23182_ (.A(_07544_),
    .B(net184),
    .C(_13198_),
    .X(_13199_));
 sky130_fd_sc_hd__a2bb2oi_2 _23183_ (.A1_N(net340),
    .A2_N(_04184_),
    .B1(_13193_),
    .B2(_13197_),
    .Y(_13200_));
 sky130_fd_sc_hd__o211ai_4 _23184_ (.A1(net341),
    .A2(_04184_),
    .B1(_13181_),
    .C1(_13192_),
    .Y(_13201_));
 sky130_fd_sc_hd__o311a_2 _23185_ (.A1(_07227_),
    .A2(_07229_),
    .A3(_13179_),
    .B1(_04227_),
    .C1(_13197_),
    .X(_13202_));
 sky130_fd_sc_hd__o211ai_4 _23186_ (.A1(net185),
    .A2(_13179_),
    .B1(_04227_),
    .C1(_13197_),
    .Y(_13203_));
 sky130_fd_sc_hd__a22oi_1 _23187_ (.A1(_02148_),
    .A2(_12718_),
    .B1(_12727_),
    .B2(_12729_),
    .Y(_13204_));
 sky130_fd_sc_hd__o2bb2ai_1 _23188_ (.A1_N(_12727_),
    .A2_N(_12729_),
    .B1(_02137_),
    .B2(_12719_),
    .Y(_13205_));
 sky130_fd_sc_hd__a31oi_2 _23189_ (.A1(_12723_),
    .A2(_12727_),
    .A3(_12729_),
    .B1(_12720_),
    .Y(_13206_));
 sky130_fd_sc_hd__o2111ai_1 _23190_ (.A1(_12722_),
    .A2(_12730_),
    .B1(_13201_),
    .C1(_13203_),
    .D1(_12721_),
    .Y(_13208_));
 sky130_fd_sc_hd__o22ai_1 _23191_ (.A1(_12720_),
    .A2(_12733_),
    .B1(_13200_),
    .B2(_13202_),
    .Y(_13209_));
 sky130_fd_sc_hd__nand3_2 _23192_ (.A(_13209_),
    .B(net163),
    .C(_13208_),
    .Y(_13210_));
 sky130_fd_sc_hd__a211o_1 _23193_ (.A1(_13193_),
    .A2(_13197_),
    .B1(_07544_),
    .C1(net184),
    .X(_13211_));
 sky130_fd_sc_hd__o2bb2ai_1 _23194_ (.A1_N(_13201_),
    .A2_N(_13203_),
    .B1(_13204_),
    .B2(_12722_),
    .Y(_13212_));
 sky130_fd_sc_hd__o2111ai_1 _23195_ (.A1(_12718_),
    .A2(_02148_),
    .B1(_13203_),
    .C1(_13201_),
    .D1(_13205_),
    .Y(_13213_));
 sky130_fd_sc_hd__nand3_2 _23196_ (.A(_13212_),
    .B(_13213_),
    .C(net163),
    .Y(_13214_));
 sky130_fd_sc_hd__o21ai_4 _23197_ (.A1(net163),
    .A2(_13198_),
    .B1(_13210_),
    .Y(_13215_));
 sky130_fd_sc_hd__o21ai_2 _23198_ (.A1(_07909_),
    .A2(_07911_),
    .B1(_13215_),
    .Y(_13216_));
 sky130_fd_sc_hd__a2bb2oi_1 _23199_ (.A1_N(_02049_),
    .A2_N(net343),
    .B1(_13211_),
    .B2(_13214_),
    .Y(_13217_));
 sky130_fd_sc_hd__o211ai_4 _23200_ (.A1(_02049_),
    .A2(net343),
    .B1(_13199_),
    .C1(_13210_),
    .Y(_13219_));
 sky130_fd_sc_hd__o211a_1 _23201_ (.A1(_02093_),
    .A2(_02115_),
    .B1(_13211_),
    .C1(_13214_),
    .X(_13220_));
 sky130_fd_sc_hd__o211ai_4 _23202_ (.A1(_02093_),
    .A2(_02115_),
    .B1(_13211_),
    .C1(_13214_),
    .Y(_13221_));
 sky130_fd_sc_hd__o21a_2 _23203_ (.A1(_00240_),
    .A2(_12738_),
    .B1(_12748_),
    .X(_13222_));
 sky130_fd_sc_hd__o21ai_2 _23204_ (.A1(_00240_),
    .A2(_12738_),
    .B1(_12748_),
    .Y(_13223_));
 sky130_fd_sc_hd__o22a_1 _23205_ (.A1(_12741_),
    .A2(_12736_),
    .B1(_12747_),
    .B2(_12744_),
    .X(_13224_));
 sky130_fd_sc_hd__nand4_4 _23206_ (.A(_12743_),
    .B(_13219_),
    .C(_13221_),
    .D(_13223_),
    .Y(_13225_));
 sky130_fd_sc_hd__o2bb2ai_4 _23207_ (.A1_N(_13219_),
    .A2_N(_13221_),
    .B1(_13222_),
    .B2(_12742_),
    .Y(_13226_));
 sky130_fd_sc_hd__o211ai_2 _23208_ (.A1(_12742_),
    .A2(_13222_),
    .B1(_13221_),
    .C1(_13219_),
    .Y(_13227_));
 sky130_fd_sc_hd__o21ai_1 _23209_ (.A1(_13217_),
    .A2(_13220_),
    .B1(_13224_),
    .Y(_13228_));
 sky130_fd_sc_hd__o211ai_4 _23210_ (.A1(_07912_),
    .A2(_07914_),
    .B1(_13227_),
    .C1(_13228_),
    .Y(_13230_));
 sky130_fd_sc_hd__and3_2 _23211_ (.A(_07917_),
    .B(_13199_),
    .C(_13210_),
    .X(_13231_));
 sky130_fd_sc_hd__nand3_1 _23212_ (.A(_13226_),
    .B(net161),
    .C(_13225_),
    .Y(_13232_));
 sky130_fd_sc_hd__a31oi_4 _23213_ (.A1(_13226_),
    .A2(net161),
    .A3(_13225_),
    .B1(_13231_),
    .Y(_13233_));
 sky130_fd_sc_hd__inv_2 _23214_ (.A(_13233_),
    .Y(_13234_));
 sky130_fd_sc_hd__and3_1 _23215_ (.A(_08301_),
    .B(_13216_),
    .C(_13230_),
    .X(_13235_));
 sky130_fd_sc_hd__or3_1 _23216_ (.A(net180),
    .B(_08298_),
    .C(_13233_),
    .X(_13236_));
 sky130_fd_sc_hd__a311oi_4 _23217_ (.A1(_13226_),
    .A2(net161),
    .A3(_13225_),
    .B1(_13231_),
    .C1(_00251_),
    .Y(_13237_));
 sky130_fd_sc_hd__o2111ai_4 _23218_ (.A1(_13215_),
    .A2(net161),
    .B1(_00207_),
    .C1(_00185_),
    .D1(_13232_),
    .Y(_13238_));
 sky130_fd_sc_hd__o211a_1 _23219_ (.A1(_00174_),
    .A2(net344),
    .B1(_13216_),
    .C1(_13230_),
    .X(_13239_));
 sky130_fd_sc_hd__o211ai_4 _23220_ (.A1(_00174_),
    .A2(net344),
    .B1(_13216_),
    .C1(_13230_),
    .Y(_13241_));
 sky130_fd_sc_hd__a21oi_1 _23221_ (.A1(_12899_),
    .A2(_12756_),
    .B1(_12760_),
    .Y(_13242_));
 sky130_fd_sc_hd__o21ai_1 _23222_ (.A1(_12325_),
    .A2(_12758_),
    .B1(_12765_),
    .Y(_13243_));
 sky130_fd_sc_hd__nand2_1 _23223_ (.A(_12763_),
    .B(_12760_),
    .Y(_13244_));
 sky130_fd_sc_hd__a21oi_2 _23224_ (.A1(_12763_),
    .A2(_12760_),
    .B1(_12764_),
    .Y(_13245_));
 sky130_fd_sc_hd__o2bb2ai_2 _23225_ (.A1_N(_13238_),
    .A2_N(_13241_),
    .B1(_13242_),
    .B2(_12762_),
    .Y(_13246_));
 sky130_fd_sc_hd__a2bb2oi_1 _23226_ (.A1_N(_00240_),
    .A2_N(_13233_),
    .B1(_13244_),
    .B2(_12765_),
    .Y(_13247_));
 sky130_fd_sc_hd__o2111ai_4 _23227_ (.A1(_12899_),
    .A2(_12756_),
    .B1(_13238_),
    .C1(_13241_),
    .D1(_13243_),
    .Y(_13248_));
 sky130_fd_sc_hd__o311a_1 _23228_ (.A1(_13237_),
    .A2(_13245_),
    .A3(_13239_),
    .B1(_08300_),
    .C1(_13246_),
    .X(_13249_));
 sky130_fd_sc_hd__o211ai_2 _23229_ (.A1(net180),
    .A2(_08298_),
    .B1(_13246_),
    .C1(_13248_),
    .Y(_13250_));
 sky130_fd_sc_hd__a31o_2 _23230_ (.A1(_13246_),
    .A2(_13248_),
    .A3(_08300_),
    .B1(_13235_),
    .X(_13252_));
 sky130_fd_sc_hd__inv_2 _23231_ (.A(_13252_),
    .Y(_13253_));
 sky130_fd_sc_hd__a21oi_1 _23232_ (.A1(_12775_),
    .A2(_11309_),
    .B1(_12785_),
    .Y(_13254_));
 sky130_fd_sc_hd__a21oi_1 _23233_ (.A1(_12776_),
    .A2(_11298_),
    .B1(_12784_),
    .Y(_13255_));
 sky130_fd_sc_hd__a32oi_2 _23234_ (.A1(_11298_),
    .A2(_12771_),
    .A3(_12774_),
    .B1(_12780_),
    .B2(_12784_),
    .Y(_13256_));
 sky130_fd_sc_hd__a311oi_4 _23235_ (.A1(_13246_),
    .A2(_13248_),
    .A3(_08300_),
    .B1(_13235_),
    .C1(_12899_),
    .Y(_13257_));
 sky130_fd_sc_hd__o221ai_2 _23236_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_08300_),
    .B2(_13233_),
    .C1(_13250_),
    .Y(_13258_));
 sky130_fd_sc_hd__a2bb2oi_1 _23237_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_13236_),
    .B2(_13250_),
    .Y(_13259_));
 sky130_fd_sc_hd__o22ai_2 _23238_ (.A1(net361),
    .A2(net345),
    .B1(_13235_),
    .B2(_13249_),
    .Y(_13260_));
 sky130_fd_sc_hd__o211ai_1 _23239_ (.A1(_12781_),
    .A2(_13254_),
    .B1(_13258_),
    .C1(_13260_),
    .Y(_13261_));
 sky130_fd_sc_hd__o22ai_1 _23240_ (.A1(_12778_),
    .A2(_13255_),
    .B1(_13257_),
    .B2(_13259_),
    .Y(_13263_));
 sky130_fd_sc_hd__nand3_1 _23241_ (.A(_13261_),
    .B(_13263_),
    .C(_08714_),
    .Y(_13264_));
 sky130_fd_sc_hd__a22o_1 _23242_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_13236_),
    .B2(_13250_),
    .X(_13265_));
 sky130_fd_sc_hd__nand3_1 _23243_ (.A(_13260_),
    .B(_13256_),
    .C(_13258_),
    .Y(_13266_));
 sky130_fd_sc_hd__o22ai_1 _23244_ (.A1(_12781_),
    .A2(_13254_),
    .B1(_13257_),
    .B2(_13259_),
    .Y(_13267_));
 sky130_fd_sc_hd__o211ai_2 _23245_ (.A1(net158),
    .A2(_08712_),
    .B1(_13266_),
    .C1(_13267_),
    .Y(_13268_));
 sky130_fd_sc_hd__o31a_2 _23246_ (.A1(net158),
    .A2(_08712_),
    .A3(_13253_),
    .B1(_13268_),
    .X(_13269_));
 sky130_fd_sc_hd__inv_2 _23247_ (.A(_13269_),
    .Y(_13270_));
 sky130_fd_sc_hd__o211ai_4 _23248_ (.A1(_13252_),
    .A2(_08714_),
    .B1(_11309_),
    .C1(_13264_),
    .Y(_13271_));
 sky130_fd_sc_hd__o211a_2 _23249_ (.A1(_08714_),
    .A2(_13253_),
    .B1(_11298_),
    .C1(_13268_),
    .X(_13272_));
 sky130_fd_sc_hd__nand3_2 _23250_ (.A(_13268_),
    .B(_11298_),
    .C(_13265_),
    .Y(_13274_));
 sky130_fd_sc_hd__o31a_1 _23251_ (.A1(_10015_),
    .A2(_12777_),
    .A3(_12788_),
    .B1(_12797_),
    .X(_13275_));
 sky130_fd_sc_hd__a21oi_1 _23252_ (.A1(_12795_),
    .A2(_12798_),
    .B1(_12792_),
    .Y(_13276_));
 sky130_fd_sc_hd__o2111ai_1 _23253_ (.A1(_12794_),
    .A2(_12797_),
    .B1(_13271_),
    .C1(_13274_),
    .D1(_12793_),
    .Y(_13277_));
 sky130_fd_sc_hd__a22o_1 _23254_ (.A1(_12793_),
    .A2(_12802_),
    .B1(_13271_),
    .B2(_13274_),
    .X(_13278_));
 sky130_fd_sc_hd__o211ai_2 _23255_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_13277_),
    .C1(_13278_),
    .Y(_13279_));
 sky130_fd_sc_hd__or3_1 _23256_ (.A(_09120_),
    .B(_09121_),
    .C(_13269_),
    .X(_13280_));
 sky130_fd_sc_hd__o2bb2ai_1 _23257_ (.A1_N(_13271_),
    .A2_N(_13274_),
    .B1(_13275_),
    .B2(_12794_),
    .Y(_13281_));
 sky130_fd_sc_hd__o21ai_1 _23258_ (.A1(_12792_),
    .A2(_12800_),
    .B1(_13271_),
    .Y(_13282_));
 sky130_fd_sc_hd__o221ai_4 _23259_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_13272_),
    .B2(_13282_),
    .C1(_13281_),
    .Y(_13283_));
 sky130_fd_sc_hd__o21ai_4 _23260_ (.A1(_09125_),
    .A2(_13269_),
    .B1(_13283_),
    .Y(_13285_));
 sky130_fd_sc_hd__or3_1 _23261_ (.A(_09553_),
    .B(net155),
    .C(_13285_),
    .X(_13286_));
 sky130_fd_sc_hd__o211ai_4 _23262_ (.A1(_13270_),
    .A2(_09125_),
    .B1(_10025_),
    .C1(_13279_),
    .Y(_13287_));
 sky130_fd_sc_hd__o221ai_4 _23263_ (.A1(net365),
    .A2(net362),
    .B1(_09125_),
    .B2(_13269_),
    .C1(_13283_),
    .Y(_13288_));
 sky130_fd_sc_hd__nand2_1 _23264_ (.A(_13287_),
    .B(_13288_),
    .Y(_13289_));
 sky130_fd_sc_hd__a32oi_2 _23265_ (.A1(_12803_),
    .A2(_12804_),
    .A3(_08907_),
    .B1(_12369_),
    .B2(_12381_),
    .Y(_13290_));
 sky130_fd_sc_hd__a21oi_2 _23266_ (.A1(_12808_),
    .A2(_12810_),
    .B1(_12811_),
    .Y(_13291_));
 sky130_fd_sc_hd__o2111ai_4 _23267_ (.A1(_12807_),
    .A2(_12809_),
    .B1(_12813_),
    .C1(_13287_),
    .D1(_13288_),
    .Y(_13292_));
 sky130_fd_sc_hd__o2bb2ai_1 _23268_ (.A1_N(_13287_),
    .A2_N(_13288_),
    .B1(_13290_),
    .B2(_12811_),
    .Y(_13293_));
 sky130_fd_sc_hd__o2111ai_4 _23269_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .C1(_13292_),
    .D1(_13293_),
    .Y(_13294_));
 sky130_fd_sc_hd__o21ai_1 _23270_ (.A1(_12811_),
    .A2(_13290_),
    .B1(_13288_),
    .Y(_13296_));
 sky130_fd_sc_hd__o21ai_4 _23271_ (.A1(net143),
    .A2(_13285_),
    .B1(_13294_),
    .Y(_13297_));
 sky130_fd_sc_hd__a21oi_1 _23272_ (.A1(_13286_),
    .A2(_13294_),
    .B1(_08918_),
    .Y(_13298_));
 sky130_fd_sc_hd__o21ai_1 _23273_ (.A1(_08863_),
    .A2(_08885_),
    .B1(_13297_),
    .Y(_13299_));
 sky130_fd_sc_hd__o211a_1 _23274_ (.A1(_13285_),
    .A2(net143),
    .B1(_08918_),
    .C1(_13294_),
    .X(_13300_));
 sky130_fd_sc_hd__o211ai_2 _23275_ (.A1(_13285_),
    .A2(net143),
    .B1(_08918_),
    .C1(_13294_),
    .Y(_13301_));
 sky130_fd_sc_hd__o211ai_2 _23276_ (.A1(_12824_),
    .A2(_12835_),
    .B1(_13299_),
    .C1(_13301_),
    .Y(_13302_));
 sky130_fd_sc_hd__o21ai_1 _23277_ (.A1(_13298_),
    .A2(_13300_),
    .B1(_12879_),
    .Y(_13303_));
 sky130_fd_sc_hd__o211ai_4 _23278_ (.A1(_09571_),
    .A2(_09573_),
    .B1(_13302_),
    .C1(_13303_),
    .Y(_13304_));
 sky130_fd_sc_hd__or3_1 _23279_ (.A(_09571_),
    .B(_09573_),
    .C(_13297_),
    .X(_13305_));
 sky130_fd_sc_hd__a21oi_2 _23280_ (.A1(_13304_),
    .A2(_13305_),
    .B1(_07888_),
    .Y(_13307_));
 sky130_fd_sc_hd__o221a_1 _23281_ (.A1(net368),
    .A2(_07866_),
    .B1(_09579_),
    .B2(_13297_),
    .C1(_13304_),
    .X(_13308_));
 sky130_fd_sc_hd__o221ai_4 _23282_ (.A1(net368),
    .A2(_07866_),
    .B1(_09579_),
    .B2(_13297_),
    .C1(_13304_),
    .Y(_13309_));
 sky130_fd_sc_hd__nand3_2 _23283_ (.A(_12395_),
    .B(_12400_),
    .C(_12841_),
    .Y(_13310_));
 sky130_fd_sc_hd__o21ai_1 _23284_ (.A1(_07044_),
    .A2(_12838_),
    .B1(_13310_),
    .Y(_13311_));
 sky130_fd_sc_hd__a211o_1 _23285_ (.A1(_13304_),
    .A2(_13305_),
    .B1(_10474_),
    .C1(net138),
    .X(_13312_));
 sky130_fd_sc_hd__o21ai_1 _23286_ (.A1(_13307_),
    .A2(_13308_),
    .B1(_13311_),
    .Y(_13313_));
 sky130_fd_sc_hd__o211ai_2 _23287_ (.A1(_07044_),
    .A2(_12838_),
    .B1(_13309_),
    .C1(_13310_),
    .Y(_13314_));
 sky130_fd_sc_hd__o211ai_4 _23288_ (.A1(_13314_),
    .A2(_13307_),
    .B1(_10480_),
    .C1(_13313_),
    .Y(_13315_));
 sky130_fd_sc_hd__nand2_1 _23289_ (.A(_13312_),
    .B(_13315_),
    .Y(_13316_));
 sky130_fd_sc_hd__o211ai_2 _23290_ (.A1(_06989_),
    .A2(net375),
    .B1(_13312_),
    .C1(_13315_),
    .Y(_13318_));
 sky130_fd_sc_hd__a22o_1 _23291_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_13312_),
    .B2(_13315_),
    .X(_13319_));
 sky130_fd_sc_hd__o2111a_1 _23292_ (.A1(_12849_),
    .A2(_06332_),
    .B1(_13318_),
    .C1(_12858_),
    .D1(_13319_),
    .X(_13320_));
 sky130_fd_sc_hd__a22oi_1 _23293_ (.A1(_12851_),
    .A2(_12858_),
    .B1(_13318_),
    .B2(_13319_),
    .Y(_13321_));
 sky130_fd_sc_hd__o21ai_1 _23294_ (.A1(_13320_),
    .A2(_13321_),
    .B1(_10954_),
    .Y(_13322_));
 sky130_fd_sc_hd__a211o_1 _23295_ (.A1(_13312_),
    .A2(_13315_),
    .B1(_10949_),
    .C1(net136),
    .X(_13323_));
 sky130_fd_sc_hd__and2_1 _23296_ (.A(_13322_),
    .B(_13323_),
    .X(_13324_));
 sky130_fd_sc_hd__or3_1 _23297_ (.A(net381),
    .B(_06310_),
    .C(_13324_),
    .X(_13325_));
 sky130_fd_sc_hd__o21ai_1 _23298_ (.A1(net381),
    .A2(_06310_),
    .B1(_13324_),
    .Y(_13326_));
 sky130_fd_sc_hd__a31o_1 _23299_ (.A1(_12859_),
    .A2(_12860_),
    .A3(_12863_),
    .B1(_12862_),
    .X(_13327_));
 sky130_fd_sc_hd__inv_2 _23300_ (.A(_13327_),
    .Y(_13329_));
 sky130_fd_sc_hd__a21oi_1 _23301_ (.A1(_13325_),
    .A2(_13326_),
    .B1(_13329_),
    .Y(_13330_));
 sky130_fd_sc_hd__a31o_1 _23302_ (.A1(_06332_),
    .A2(_13322_),
    .A3(_13323_),
    .B1(_13327_),
    .X(_13331_));
 sky130_fd_sc_hd__and3_1 _23303_ (.A(_13325_),
    .B(_13326_),
    .C(_13329_),
    .X(_13332_));
 sky130_fd_sc_hd__or3_1 _23304_ (.A(_11459_),
    .B(_11461_),
    .C(_13324_),
    .X(_13333_));
 sky130_fd_sc_hd__o31ai_2 _23305_ (.A1(_11464_),
    .A2(_13330_),
    .A3(_13332_),
    .B1(_13333_),
    .Y(_13334_));
 sky130_fd_sc_hd__a21oi_1 _23306_ (.A1(_12870_),
    .A2(_12872_),
    .B1(_12873_),
    .Y(_13335_));
 sky130_fd_sc_hd__a211o_1 _23307_ (.A1(_12870_),
    .A2(_12872_),
    .B1(_12873_),
    .C1(_05862_),
    .X(_13336_));
 sky130_fd_sc_hd__a21oi_1 _23308_ (.A1(net395),
    .A2(_05796_),
    .B1(_13335_),
    .Y(_13337_));
 sky130_fd_sc_hd__a21oi_2 _23309_ (.A1(_11943_),
    .A2(_13336_),
    .B1(_13334_),
    .Y(_13338_));
 sky130_fd_sc_hd__xnor2_1 _23310_ (.A(_12878_),
    .B(_13338_),
    .Y(net92));
 sky130_fd_sc_hd__o2111ai_4 _23311_ (.A1(_11944_),
    .A2(_12871_),
    .B1(_12868_),
    .C1(_12418_),
    .D1(_13338_),
    .Y(_13340_));
 sky130_fd_sc_hd__o211a_2 _23312_ (.A1(_12880_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_12887_),
    .X(_13341_));
 sky130_fd_sc_hd__o311a_1 _23313_ (.A1(_11470_),
    .A2(_12882_),
    .A3(_12886_),
    .B1(_07724_),
    .C1(net357),
    .X(_13342_));
 sky130_fd_sc_hd__or4_2 _23314_ (.A(_06848_),
    .B(net374),
    .C(_07702_),
    .D(_13341_),
    .X(_13343_));
 sky130_fd_sc_hd__o311a_1 _23315_ (.A1(_11470_),
    .A2(_12882_),
    .A3(_12886_),
    .B1(_10971_),
    .C1(net357),
    .X(_13344_));
 sky130_fd_sc_hd__o22a_1 _23316_ (.A1(_10965_),
    .A2(_10967_),
    .B1(_06848_),
    .B2(_13341_),
    .X(_13345_));
 sky130_fd_sc_hd__nor2_1 _23317_ (.A(_13344_),
    .B(_13345_),
    .Y(_13346_));
 sky130_fd_sc_hd__o32ai_4 _23318_ (.A1(net150),
    .A2(_12891_),
    .A3(_12892_),
    .B1(_12898_),
    .B2(_12900_),
    .Y(_13347_));
 sky130_fd_sc_hd__nand2_2 _23319_ (.A(_13347_),
    .B(_13346_),
    .Y(_13348_));
 sky130_fd_sc_hd__o221ai_4 _23320_ (.A1(_13344_),
    .A2(_13345_),
    .B1(_12898_),
    .B2(_12900_),
    .C1(_12896_),
    .Y(_13350_));
 sky130_fd_sc_hd__o221ai_4 _23321_ (.A1(net374),
    .A2(_07702_),
    .B1(_13346_),
    .B2(_13347_),
    .C1(_13348_),
    .Y(_13351_));
 sky130_fd_sc_hd__a31oi_2 _23322_ (.A1(_13348_),
    .A2(_13350_),
    .A3(net355),
    .B1(_13342_),
    .Y(_13352_));
 sky130_fd_sc_hd__a21oi_2 _23323_ (.A1(_13343_),
    .A2(_13351_),
    .B1(net338),
    .Y(_13353_));
 sky130_fd_sc_hd__or3_1 _23324_ (.A(_08678_),
    .B(_08700_),
    .C(_13352_),
    .X(_13354_));
 sky130_fd_sc_hd__a2bb2oi_2 _23325_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_13343_),
    .B2(_13351_),
    .Y(_13355_));
 sky130_fd_sc_hd__or3_1 _23326_ (.A(_10489_),
    .B(_10490_),
    .C(_13352_),
    .X(_13356_));
 sky130_fd_sc_hd__a31oi_1 _23327_ (.A1(_13348_),
    .A2(_13350_),
    .A3(net355),
    .B1(_10492_),
    .Y(_13357_));
 sky130_fd_sc_hd__o311a_2 _23328_ (.A1(_06848_),
    .A2(net355),
    .A3(_13341_),
    .B1(net150),
    .C1(_13351_),
    .X(_13358_));
 sky130_fd_sc_hd__a21oi_1 _23329_ (.A1(_13343_),
    .A2(_13357_),
    .B1(_13355_),
    .Y(_13359_));
 sky130_fd_sc_hd__a31oi_2 _23330_ (.A1(_12913_),
    .A2(_12918_),
    .A3(_12922_),
    .B1(_12909_),
    .Y(_13361_));
 sky130_fd_sc_hd__a31o_1 _23331_ (.A1(_12913_),
    .A2(_12918_),
    .A3(_12922_),
    .B1(_12909_),
    .X(_13362_));
 sky130_fd_sc_hd__o221ai_4 _23332_ (.A1(_10026_),
    .A2(_12906_),
    .B1(_13355_),
    .B2(_13358_),
    .C1(_12926_),
    .Y(_13363_));
 sky130_fd_sc_hd__nand2_2 _23333_ (.A(_13362_),
    .B(_13359_),
    .Y(_13364_));
 sky130_fd_sc_hd__o211ai_2 _23334_ (.A1(_08678_),
    .A2(_08700_),
    .B1(_13363_),
    .C1(_13364_),
    .Y(_13365_));
 sky130_fd_sc_hd__o31a_2 _23335_ (.A1(_08678_),
    .A2(_08700_),
    .A3(_13352_),
    .B1(_13365_),
    .X(_13366_));
 sky130_fd_sc_hd__a21oi_1 _23336_ (.A1(_13354_),
    .A2(_13365_),
    .B1(net335),
    .Y(_13367_));
 sky130_fd_sc_hd__or3_1 _23337_ (.A(net351),
    .B(_09807_),
    .C(_13366_),
    .X(_13368_));
 sky130_fd_sc_hd__a2bb2oi_2 _23338_ (.A1_N(net170),
    .A2_N(net169),
    .B1(_13354_),
    .B2(_13365_),
    .Y(_13369_));
 sky130_fd_sc_hd__a2bb2o_1 _23339_ (.A1_N(net170),
    .A2_N(net169),
    .B1(_13354_),
    .B2(_13365_),
    .X(_13370_));
 sky130_fd_sc_hd__a311oi_4 _23340_ (.A1(_13364_),
    .A2(net338),
    .A3(_13363_),
    .B1(net151),
    .C1(_13353_),
    .Y(_13372_));
 sky130_fd_sc_hd__a311o_1 _23341_ (.A1(_13364_),
    .A2(net338),
    .A3(_13363_),
    .B1(net151),
    .C1(_13353_),
    .X(_13373_));
 sky130_fd_sc_hd__nand3_2 _23342_ (.A(_12042_),
    .B(_12045_),
    .C(_11568_),
    .Y(_13374_));
 sky130_fd_sc_hd__a21oi_1 _23343_ (.A1(net173),
    .A2(_12481_),
    .B1(_13374_),
    .Y(_13375_));
 sky130_fd_sc_hd__o21bai_4 _23344_ (.A1(_13375_),
    .A2(_12934_),
    .B1_N(_12484_),
    .Y(_13376_));
 sky130_fd_sc_hd__o41ai_4 _23345_ (.A1(_11578_),
    .A2(_12484_),
    .A3(_13374_),
    .A4(_12486_),
    .B1(_12946_),
    .Y(_13377_));
 sky130_fd_sc_hd__o22a_1 _23346_ (.A1(net172),
    .A2(_12933_),
    .B1(_13376_),
    .B2(_13377_),
    .X(_13378_));
 sky130_fd_sc_hd__o22ai_2 _23347_ (.A1(net172),
    .A2(_12933_),
    .B1(_13376_),
    .B2(_13377_),
    .Y(_13379_));
 sky130_fd_sc_hd__o221ai_4 _23348_ (.A1(_13377_),
    .A2(_13376_),
    .B1(_13372_),
    .B2(_13369_),
    .C1(_12944_),
    .Y(_13380_));
 sky130_fd_sc_hd__nand3_2 _23349_ (.A(_13370_),
    .B(_13373_),
    .C(_13379_),
    .Y(_13381_));
 sky130_fd_sc_hd__nand3_2 _23350_ (.A(_13381_),
    .B(net335),
    .C(_13380_),
    .Y(_13383_));
 sky130_fd_sc_hd__o31a_2 _23351_ (.A1(net351),
    .A2(_09807_),
    .A3(_13366_),
    .B1(_13383_),
    .X(_13384_));
 sky130_fd_sc_hd__a211o_1 _23352_ (.A1(_13368_),
    .A2(_13383_),
    .B1(_11046_),
    .C1(_11057_),
    .X(_13385_));
 sky130_fd_sc_hd__o211a_1 _23353_ (.A1(_12502_),
    .A2(_12499_),
    .B1(_12498_),
    .C1(_12951_),
    .X(_13386_));
 sky130_fd_sc_hd__o211ai_2 _23354_ (.A1(_12502_),
    .A2(_12499_),
    .B1(_12498_),
    .C1(_12951_),
    .Y(_13387_));
 sky130_fd_sc_hd__a2bb2oi_2 _23355_ (.A1_N(_09588_),
    .A2_N(_09590_),
    .B1(_13368_),
    .B2(_13383_),
    .Y(_13388_));
 sky130_fd_sc_hd__a22o_2 _23356_ (.A1(_09589_),
    .A2(_09591_),
    .B1(_13368_),
    .B2(_13383_),
    .X(_13389_));
 sky130_fd_sc_hd__a311oi_4 _23357_ (.A1(_13381_),
    .A2(net335),
    .A3(_13380_),
    .B1(_09595_),
    .C1(_13367_),
    .Y(_13390_));
 sky130_fd_sc_hd__o211ai_4 _23358_ (.A1(net335),
    .A2(_13366_),
    .B1(net172),
    .C1(_13383_),
    .Y(_13391_));
 sky130_fd_sc_hd__o211ai_4 _23359_ (.A1(net173),
    .A2(_12950_),
    .B1(_13387_),
    .C1(_13391_),
    .Y(_13392_));
 sky130_fd_sc_hd__o22ai_2 _23360_ (.A1(_12952_),
    .A2(_13386_),
    .B1(_13388_),
    .B2(_13390_),
    .Y(_13394_));
 sky130_fd_sc_hd__o211ai_4 _23361_ (.A1(_13388_),
    .A2(_13392_),
    .B1(net332),
    .C1(_13394_),
    .Y(_13395_));
 sky130_fd_sc_hd__o21ai_2 _23362_ (.A1(net332),
    .A2(_13384_),
    .B1(_13395_),
    .Y(_13396_));
 sky130_fd_sc_hd__a2bb2oi_4 _23363_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_13385_),
    .B2(_13395_),
    .Y(_13397_));
 sky130_fd_sc_hd__a2bb2o_1 _23364_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_13385_),
    .B2(_13395_),
    .X(_13398_));
 sky130_fd_sc_hd__o211a_2 _23365_ (.A1(net332),
    .A2(_13384_),
    .B1(net174),
    .C1(_13395_),
    .X(_13399_));
 sky130_fd_sc_hd__o211ai_4 _23366_ (.A1(net332),
    .A2(_13384_),
    .B1(net174),
    .C1(_13395_),
    .Y(_13400_));
 sky130_fd_sc_hd__nor2_1 _23367_ (.A(_13397_),
    .B(_13399_),
    .Y(_13401_));
 sky130_fd_sc_hd__nand3_2 _23368_ (.A(_12517_),
    .B(_12968_),
    .C(_12972_),
    .Y(_13402_));
 sky130_fd_sc_hd__o21ai_1 _23369_ (.A1(net175),
    .A2(_12964_),
    .B1(_13402_),
    .Y(_13403_));
 sky130_fd_sc_hd__nand3_1 _23370_ (.A(_13398_),
    .B(_13400_),
    .C(_13403_),
    .Y(_13405_));
 sky130_fd_sc_hd__o221ai_2 _23371_ (.A1(net175),
    .A2(_12964_),
    .B1(_13397_),
    .B2(_13399_),
    .C1(_13402_),
    .Y(_13406_));
 sky130_fd_sc_hd__o211ai_2 _23372_ (.A1(net329),
    .A2(net327),
    .B1(_13405_),
    .C1(_13406_),
    .Y(_13407_));
 sky130_fd_sc_hd__a211o_1 _23373_ (.A1(_13385_),
    .A2(_13395_),
    .B1(net329),
    .C1(net327),
    .X(_13408_));
 sky130_fd_sc_hd__o21ai_1 _23374_ (.A1(_13397_),
    .A2(_13399_),
    .B1(_13403_),
    .Y(_13409_));
 sky130_fd_sc_hd__nand4_1 _23375_ (.A(_12970_),
    .B(_13398_),
    .C(_13400_),
    .D(_13402_),
    .Y(_13410_));
 sky130_fd_sc_hd__o211ai_2 _23376_ (.A1(net329),
    .A2(net327),
    .B1(_13409_),
    .C1(_13410_),
    .Y(_13411_));
 sky130_fd_sc_hd__o21a_2 _23377_ (.A1(net311),
    .A2(_13396_),
    .B1(_13407_),
    .X(_13412_));
 sky130_fd_sc_hd__o211ai_4 _23378_ (.A1(_13396_),
    .A2(net311),
    .B1(net175),
    .C1(_13407_),
    .Y(_13413_));
 sky130_fd_sc_hd__o211ai_4 _23379_ (.A1(_08728_),
    .A2(net195),
    .B1(_13408_),
    .C1(_13411_),
    .Y(_13414_));
 sky130_fd_sc_hd__nand2_1 _23380_ (.A(_13413_),
    .B(_13414_),
    .Y(_13416_));
 sky130_fd_sc_hd__o211ai_2 _23381_ (.A1(_12992_),
    .A2(_12539_),
    .B1(_12984_),
    .C1(_12991_),
    .Y(_13417_));
 sky130_fd_sc_hd__o211ai_4 _23382_ (.A1(net199),
    .A2(_12978_),
    .B1(_12996_),
    .C1(_13416_),
    .Y(_13418_));
 sky130_fd_sc_hd__o2111ai_4 _23383_ (.A1(_12981_),
    .A2(_12994_),
    .B1(_13413_),
    .C1(_13414_),
    .D1(_12984_),
    .Y(_13419_));
 sky130_fd_sc_hd__o211ai_4 _23384_ (.A1(_00011_),
    .A2(net323),
    .B1(_13418_),
    .C1(_13419_),
    .Y(_13420_));
 sky130_fd_sc_hd__a2bb2o_2 _23385_ (.A1_N(_14458_),
    .A2_N(_00000_),
    .B1(_13408_),
    .B2(_13411_),
    .X(_13421_));
 sky130_fd_sc_hd__inv_2 _23386_ (.A(_13421_),
    .Y(_13422_));
 sky130_fd_sc_hd__a31oi_4 _23387_ (.A1(_13419_),
    .A2(net307),
    .A3(_13418_),
    .B1(_13422_),
    .Y(_13423_));
 sky130_fd_sc_hd__a31o_2 _23388_ (.A1(_13419_),
    .A2(net307),
    .A3(_13418_),
    .B1(_13422_),
    .X(_13424_));
 sky130_fd_sc_hd__a211o_2 _23389_ (.A1(_13420_),
    .A2(_13421_),
    .B1(net304),
    .C1(_01951_),
    .X(_13425_));
 sky130_fd_sc_hd__inv_2 _23390_ (.A(_13425_),
    .Y(_13427_));
 sky130_fd_sc_hd__a21oi_2 _23391_ (.A1(_13420_),
    .A2(_13421_),
    .B1(net199),
    .Y(_13428_));
 sky130_fd_sc_hd__a22o_1 _23392_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_13420_),
    .B2(_13421_),
    .X(_13429_));
 sky130_fd_sc_hd__a31o_2 _23393_ (.A1(_13419_),
    .A2(net307),
    .A3(_13418_),
    .B1(net198),
    .X(_13430_));
 sky130_fd_sc_hd__a311o_1 _23394_ (.A1(_13418_),
    .A2(_13419_),
    .A3(net307),
    .B1(_13422_),
    .C1(net198),
    .X(_13431_));
 sky130_fd_sc_hd__a41oi_2 _23395_ (.A1(_08308_),
    .A2(_08310_),
    .A3(_13420_),
    .A4(_13421_),
    .B1(_13428_),
    .Y(_13432_));
 sky130_fd_sc_hd__o21ai_1 _23396_ (.A1(_13422_),
    .A2(_13430_),
    .B1(_13429_),
    .Y(_13433_));
 sky130_fd_sc_hd__nand4_1 _23397_ (.A(_11641_),
    .B(_11644_),
    .C(_12108_),
    .D(_12111_),
    .Y(_13434_));
 sky130_fd_sc_hd__nor3_2 _23398_ (.A(_12551_),
    .B(_12552_),
    .C(_13434_),
    .Y(_13435_));
 sky130_fd_sc_hd__o21ai_1 _23399_ (.A1(_07936_),
    .A2(_13002_),
    .B1(_13435_),
    .Y(_13436_));
 sky130_fd_sc_hd__a21oi_1 _23400_ (.A1(_13006_),
    .A2(_13435_),
    .B1(_13007_),
    .Y(_13438_));
 sky130_fd_sc_hd__o211ai_4 _23401_ (.A1(_13011_),
    .A2(_13005_),
    .B1(_13008_),
    .C1(_13436_),
    .Y(_13439_));
 sky130_fd_sc_hd__o211ai_2 _23402_ (.A1(_07935_),
    .A2(_13001_),
    .B1(_13435_),
    .C1(_11659_),
    .Y(_13440_));
 sky130_fd_sc_hd__nand4_4 _23403_ (.A(_13435_),
    .B(_13008_),
    .C(_13006_),
    .D(_11659_),
    .Y(_13441_));
 sky130_fd_sc_hd__a2bb2oi_1 _23404_ (.A1_N(_13005_),
    .A2_N(_13440_),
    .B1(_13013_),
    .B2(_13438_),
    .Y(_13442_));
 sky130_fd_sc_hd__o21ai_2 _23405_ (.A1(_13005_),
    .A2(_13440_),
    .B1(_13439_),
    .Y(_13443_));
 sky130_fd_sc_hd__o211ai_1 _23406_ (.A1(_13005_),
    .A2(_13440_),
    .B1(_13439_),
    .C1(_13433_),
    .Y(_13444_));
 sky130_fd_sc_hd__nand2_1 _23407_ (.A(_13443_),
    .B(_13432_),
    .Y(_13445_));
 sky130_fd_sc_hd__nand4_2 _23408_ (.A(_13429_),
    .B(_13431_),
    .C(_13439_),
    .D(_13441_),
    .Y(_13446_));
 sky130_fd_sc_hd__a22o_1 _23409_ (.A1(_13429_),
    .A2(_13431_),
    .B1(_13439_),
    .B2(_13441_),
    .X(_13447_));
 sky130_fd_sc_hd__nand3_2 _23410_ (.A(_13447_),
    .B(net278),
    .C(_13446_),
    .Y(_13449_));
 sky130_fd_sc_hd__a311o_1 _23411_ (.A1(_13418_),
    .A2(_13419_),
    .A3(net307),
    .B1(_13422_),
    .C1(net278),
    .X(_13450_));
 sky130_fd_sc_hd__nand3_2 _23412_ (.A(_13445_),
    .B(net278),
    .C(_13444_),
    .Y(_13451_));
 sky130_fd_sc_hd__o221a_1 _23413_ (.A1(_03986_),
    .A2(_03997_),
    .B1(_13424_),
    .B2(net278),
    .C1(_13451_),
    .X(_13452_));
 sky130_fd_sc_hd__a211o_2 _23414_ (.A1(_13425_),
    .A2(_13449_),
    .B1(net302),
    .C1(_04019_),
    .X(_13453_));
 sky130_fd_sc_hd__a311oi_4 _23415_ (.A1(_13447_),
    .A2(net278),
    .A3(_13446_),
    .B1(_07936_),
    .C1(_13427_),
    .Y(_13454_));
 sky130_fd_sc_hd__nand3_4 _23416_ (.A(_13449_),
    .B(_07935_),
    .C(_13425_),
    .Y(_13455_));
 sky130_fd_sc_hd__o211ai_4 _23417_ (.A1(_13424_),
    .A2(net278),
    .B1(_07936_),
    .C1(_13451_),
    .Y(_13456_));
 sky130_fd_sc_hd__a21oi_1 _23418_ (.A1(_12564_),
    .A2(_13018_),
    .B1(_13024_),
    .Y(_13457_));
 sky130_fd_sc_hd__a31o_1 _23419_ (.A1(_12564_),
    .A2(_13018_),
    .A3(_13023_),
    .B1(_13024_),
    .X(_13458_));
 sky130_fd_sc_hd__a31oi_4 _23420_ (.A1(_12564_),
    .A2(_13018_),
    .A3(_13023_),
    .B1(_13024_),
    .Y(_13460_));
 sky130_fd_sc_hd__o2bb2ai_4 _23421_ (.A1_N(_13455_),
    .A2_N(_13456_),
    .B1(_13457_),
    .B2(_13022_),
    .Y(_13461_));
 sky130_fd_sc_hd__nand3_4 _23422_ (.A(_13458_),
    .B(_13456_),
    .C(_13455_),
    .Y(_13462_));
 sky130_fd_sc_hd__nand3_4 _23423_ (.A(_13461_),
    .B(_13462_),
    .C(net277),
    .Y(_13463_));
 sky130_fd_sc_hd__a31o_1 _23424_ (.A1(_13461_),
    .A2(_13462_),
    .A3(net277),
    .B1(_13452_),
    .X(_13464_));
 sky130_fd_sc_hd__and3_1 _23425_ (.A(_05234_),
    .B(_13453_),
    .C(_13463_),
    .X(_13465_));
 sky130_fd_sc_hd__o221ai_4 _23426_ (.A1(net227),
    .A2(_12572_),
    .B1(net224),
    .B2(_13036_),
    .C1(_13043_),
    .Y(_13466_));
 sky130_fd_sc_hd__a22oi_4 _23427_ (.A1(net224),
    .A2(_13036_),
    .B1(_13043_),
    .B2(_12576_),
    .Y(_13467_));
 sky130_fd_sc_hd__nand2_1 _23428_ (.A(_13039_),
    .B(_13466_),
    .Y(_13468_));
 sky130_fd_sc_hd__a311oi_4 _23429_ (.A1(_13461_),
    .A2(_13462_),
    .A3(net277),
    .B1(net202),
    .C1(_13452_),
    .Y(_13469_));
 sky130_fd_sc_hd__nand3_4 _23430_ (.A(_13463_),
    .B(_07564_),
    .C(_13453_),
    .Y(_13471_));
 sky130_fd_sc_hd__a2bb2oi_4 _23431_ (.A1_N(net221),
    .A2_N(_07557_),
    .B1(_13453_),
    .B2(_13463_),
    .Y(_13472_));
 sky130_fd_sc_hd__o21ai_1 _23432_ (.A1(net221),
    .A2(_07557_),
    .B1(_13464_),
    .Y(_13473_));
 sky130_fd_sc_hd__nor2_1 _23433_ (.A(_13469_),
    .B(_13472_),
    .Y(_13474_));
 sky130_fd_sc_hd__nand3_2 _23434_ (.A(_13468_),
    .B(_13471_),
    .C(_13473_),
    .Y(_13475_));
 sky130_fd_sc_hd__o22ai_4 _23435_ (.A1(_13037_),
    .A2(_13467_),
    .B1(_13469_),
    .B2(_13472_),
    .Y(_13476_));
 sky130_fd_sc_hd__o211ai_2 _23436_ (.A1(net296),
    .A2(_05232_),
    .B1(_13475_),
    .C1(_13476_),
    .Y(_13477_));
 sky130_fd_sc_hd__a21oi_1 _23437_ (.A1(_13453_),
    .A2(_13463_),
    .B1(net272),
    .Y(_13478_));
 sky130_fd_sc_hd__o211ai_2 _23438_ (.A1(_13037_),
    .A2(_13467_),
    .B1(_13471_),
    .C1(_13473_),
    .Y(_13479_));
 sky130_fd_sc_hd__o21ai_2 _23439_ (.A1(_13469_),
    .A2(_13472_),
    .B1(_13468_),
    .Y(_13480_));
 sky130_fd_sc_hd__o211ai_2 _23440_ (.A1(net296),
    .A2(_05232_),
    .B1(_13479_),
    .C1(_13480_),
    .Y(_13482_));
 sky130_fd_sc_hd__a31o_2 _23441_ (.A1(_13479_),
    .A2(_13480_),
    .A3(net272),
    .B1(_13478_),
    .X(_13483_));
 sky130_fd_sc_hd__a31o_2 _23442_ (.A1(_13475_),
    .A2(_13476_),
    .A3(net272),
    .B1(_13465_),
    .X(_13484_));
 sky130_fd_sc_hd__a311oi_2 _23443_ (.A1(_13475_),
    .A2(_13476_),
    .A3(net272),
    .B1(net224),
    .C1(_13465_),
    .Y(_13485_));
 sky130_fd_sc_hd__o211ai_4 _23444_ (.A1(_13464_),
    .A2(net272),
    .B1(net222),
    .C1(_13477_),
    .Y(_13486_));
 sky130_fd_sc_hd__a311oi_2 _23445_ (.A1(_13479_),
    .A2(_13480_),
    .A3(net272),
    .B1(net222),
    .C1(_13478_),
    .Y(_13487_));
 sky130_fd_sc_hd__nand3b_4 _23446_ (.A_N(_13478_),
    .B(_13482_),
    .C(net224),
    .Y(_13488_));
 sky130_fd_sc_hd__nand2_1 _23447_ (.A(_13486_),
    .B(_13488_),
    .Y(_13489_));
 sky130_fd_sc_hd__o21ai_2 _23448_ (.A1(net225),
    .A2(_13054_),
    .B1(_13072_),
    .Y(_13490_));
 sky130_fd_sc_hd__o22ai_2 _23449_ (.A1(net227),
    .A2(_13052_),
    .B1(_13490_),
    .B2(_13068_),
    .Y(_13491_));
 sky130_fd_sc_hd__a31oi_2 _23450_ (.A1(_13059_),
    .A2(_13069_),
    .A3(_13072_),
    .B1(_13055_),
    .Y(_13493_));
 sky130_fd_sc_hd__nand3_2 _23451_ (.A(_13491_),
    .B(_13488_),
    .C(_13486_),
    .Y(_13494_));
 sky130_fd_sc_hd__o211a_1 _23452_ (.A1(_13485_),
    .A2(_13487_),
    .B1(_13056_),
    .C1(_13080_),
    .X(_13495_));
 sky130_fd_sc_hd__o211ai_2 _23453_ (.A1(_13485_),
    .A2(_13487_),
    .B1(_13056_),
    .C1(_13080_),
    .Y(_13496_));
 sky130_fd_sc_hd__o22ai_4 _23454_ (.A1(net270),
    .A2(net268),
    .B1(_13489_),
    .B2(_13493_),
    .Y(_13497_));
 sky130_fd_sc_hd__nand3_1 _23455_ (.A(_13494_),
    .B(_13496_),
    .C(net245),
    .Y(_13498_));
 sky130_fd_sc_hd__and3_4 _23456_ (.A(_13483_),
    .B(_05484_),
    .C(_05482_),
    .X(_13499_));
 sky130_fd_sc_hd__a311o_2 _23457_ (.A1(_13475_),
    .A2(_13476_),
    .A3(net272),
    .B1(net245),
    .C1(_13465_),
    .X(_13500_));
 sky130_fd_sc_hd__o32a_4 _23458_ (.A1(net270),
    .A2(net268),
    .A3(_13484_),
    .B1(_13495_),
    .B2(_13497_),
    .X(_13501_));
 sky130_fd_sc_hd__o22ai_4 _23459_ (.A1(net245),
    .A2(_13484_),
    .B1(_13495_),
    .B2(_13497_),
    .Y(_13502_));
 sky130_fd_sc_hd__a21oi_2 _23460_ (.A1(_13498_),
    .A2(_13500_),
    .B1(net227),
    .Y(_13504_));
 sky130_fd_sc_hd__o21ai_4 _23461_ (.A1(_06914_),
    .A2(net250),
    .B1(_13502_),
    .Y(_13505_));
 sky130_fd_sc_hd__o22a_1 _23462_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_13495_),
    .B2(_13497_),
    .X(_13506_));
 sky130_fd_sc_hd__a31o_2 _23463_ (.A1(_13494_),
    .A2(_13496_),
    .A3(net245),
    .B1(net225),
    .X(_13507_));
 sky130_fd_sc_hd__a311oi_2 _23464_ (.A1(_13494_),
    .A2(_13496_),
    .A3(net245),
    .B1(_13499_),
    .C1(net225),
    .Y(_13508_));
 sky130_fd_sc_hd__a311o_1 _23465_ (.A1(_13494_),
    .A2(_13496_),
    .A3(net245),
    .B1(_13499_),
    .C1(net225),
    .X(_13509_));
 sky130_fd_sc_hd__a21oi_2 _23466_ (.A1(_13500_),
    .A2(_13506_),
    .B1(_13504_),
    .Y(_13510_));
 sky130_fd_sc_hd__o21ai_1 _23467_ (.A1(_13499_),
    .A2(_13507_),
    .B1(_13505_),
    .Y(_13511_));
 sky130_fd_sc_hd__o2111ai_4 _23468_ (.A1(_11720_),
    .A2(_11714_),
    .B1(_11719_),
    .C1(_12183_),
    .D1(_12186_),
    .Y(_13512_));
 sky130_fd_sc_hd__a211oi_4 _23469_ (.A1(_12603_),
    .A2(_12620_),
    .B1(_13512_),
    .C1(_12623_),
    .Y(_13513_));
 sky130_fd_sc_hd__nand2_1 _23470_ (.A(_13088_),
    .B(_13513_),
    .Y(_13515_));
 sky130_fd_sc_hd__a21oi_1 _23471_ (.A1(_13088_),
    .A2(_13513_),
    .B1(_13089_),
    .Y(_13516_));
 sky130_fd_sc_hd__o211ai_4 _23472_ (.A1(_13094_),
    .A2(_13087_),
    .B1(_13090_),
    .C1(_13515_),
    .Y(_13517_));
 sky130_fd_sc_hd__nand3_2 _23473_ (.A(_11725_),
    .B(_13090_),
    .C(_13513_),
    .Y(_13518_));
 sky130_fd_sc_hd__nand4_4 _23474_ (.A(_13513_),
    .B(_13090_),
    .C(_13088_),
    .D(_11725_),
    .Y(_13519_));
 sky130_fd_sc_hd__a2bb2oi_4 _23475_ (.A1_N(_13087_),
    .A2_N(_13518_),
    .B1(_13099_),
    .B2(_13516_),
    .Y(_13520_));
 sky130_fd_sc_hd__o21ai_2 _23476_ (.A1(_13087_),
    .A2(_13518_),
    .B1(_13517_),
    .Y(_13521_));
 sky130_fd_sc_hd__a21oi_2 _23477_ (.A1(_13517_),
    .A2(_13519_),
    .B1(_13511_),
    .Y(_13522_));
 sky130_fd_sc_hd__o221ai_2 _23478_ (.A1(_13087_),
    .A2(_13518_),
    .B1(_13508_),
    .B2(_13504_),
    .C1(_13517_),
    .Y(_13523_));
 sky130_fd_sc_hd__o21ai_2 _23479_ (.A1(_05750_),
    .A2(net264),
    .B1(_13523_),
    .Y(_13524_));
 sky130_fd_sc_hd__nand4_4 _23480_ (.A(_13505_),
    .B(_13509_),
    .C(_13517_),
    .D(_13519_),
    .Y(_13526_));
 sky130_fd_sc_hd__a22o_1 _23481_ (.A1(_13505_),
    .A2(_13509_),
    .B1(_13517_),
    .B2(_13519_),
    .X(_13527_));
 sky130_fd_sc_hd__a21oi_2 _23482_ (.A1(_13498_),
    .A2(_13500_),
    .B1(net243),
    .Y(_13528_));
 sky130_fd_sc_hd__or3_1 _23483_ (.A(_05750_),
    .B(net264),
    .C(_13501_),
    .X(_13529_));
 sky130_fd_sc_hd__o221ai_4 _23484_ (.A1(_05750_),
    .A2(net264),
    .B1(_13510_),
    .B2(_13520_),
    .C1(_13526_),
    .Y(_13530_));
 sky130_fd_sc_hd__a31o_1 _23485_ (.A1(_13527_),
    .A2(net243),
    .A3(_13526_),
    .B1(_13528_),
    .X(_13531_));
 sky130_fd_sc_hd__o221a_1 _23486_ (.A1(net243),
    .A2(_13502_),
    .B1(_13522_),
    .B2(_13524_),
    .C1(_05995_),
    .X(_13532_));
 sky130_fd_sc_hd__a211o_1 _23487_ (.A1(_13529_),
    .A2(_13530_),
    .B1(net260),
    .C1(net258),
    .X(_13533_));
 sky130_fd_sc_hd__a311oi_4 _23488_ (.A1(_13527_),
    .A2(net243),
    .A3(_13526_),
    .B1(_13528_),
    .C1(net232),
    .Y(_13534_));
 sky130_fd_sc_hd__nand3_4 _23489_ (.A(_13530_),
    .B(net234),
    .C(_13529_),
    .Y(_13535_));
 sky130_fd_sc_hd__o221ai_4 _23490_ (.A1(net243),
    .A2(_13502_),
    .B1(_13522_),
    .B2(_13524_),
    .C1(net233),
    .Y(_13537_));
 sky130_fd_sc_hd__o221a_1 _23491_ (.A1(_12640_),
    .A2(_12636_),
    .B1(_06314_),
    .B2(_13105_),
    .C1(_12635_),
    .X(_13538_));
 sky130_fd_sc_hd__o31a_1 _23492_ (.A1(_13102_),
    .A2(net252),
    .A3(_13100_),
    .B1(_13112_),
    .X(_13539_));
 sky130_fd_sc_hd__o21ai_1 _23493_ (.A1(_13107_),
    .A2(_13113_),
    .B1(_13111_),
    .Y(_13540_));
 sky130_fd_sc_hd__a21oi_2 _23494_ (.A1(_13109_),
    .A2(_13112_),
    .B1(_13110_),
    .Y(_13541_));
 sky130_fd_sc_hd__a21oi_1 _23495_ (.A1(_13535_),
    .A2(_13537_),
    .B1(_13540_),
    .Y(_13542_));
 sky130_fd_sc_hd__o2bb2ai_4 _23496_ (.A1_N(_13535_),
    .A2_N(_13537_),
    .B1(_13538_),
    .B2(_13107_),
    .Y(_13543_));
 sky130_fd_sc_hd__o211a_1 _23497_ (.A1(_13110_),
    .A2(_13539_),
    .B1(_13537_),
    .C1(_13535_),
    .X(_13544_));
 sky130_fd_sc_hd__o211ai_4 _23498_ (.A1(_13110_),
    .A2(_13539_),
    .B1(_13537_),
    .C1(_13535_),
    .Y(_13545_));
 sky130_fd_sc_hd__a31oi_2 _23499_ (.A1(_13535_),
    .A2(_13537_),
    .A3(_13540_),
    .B1(_05995_),
    .Y(_13546_));
 sky130_fd_sc_hd__o211ai_4 _23500_ (.A1(net260),
    .A2(net258),
    .B1(_13543_),
    .C1(_13545_),
    .Y(_13548_));
 sky130_fd_sc_hd__o22ai_2 _23501_ (.A1(net260),
    .A2(net258),
    .B1(_13542_),
    .B2(_13544_),
    .Y(_13549_));
 sky130_fd_sc_hd__a31o_2 _23502_ (.A1(net240),
    .A2(_13543_),
    .A3(_13545_),
    .B1(_13532_),
    .X(_13550_));
 sky130_fd_sc_hd__o221a_1 _23503_ (.A1(net263),
    .A2(_12650_),
    .B1(net254),
    .B2(_13124_),
    .C1(_12671_),
    .X(_13551_));
 sky130_fd_sc_hd__a31oi_4 _23504_ (.A1(_12653_),
    .A2(_12671_),
    .A3(_13127_),
    .B1(_13128_),
    .Y(_13552_));
 sky130_fd_sc_hd__a211oi_4 _23505_ (.A1(_13546_),
    .A2(_13543_),
    .B1(_13532_),
    .C1(net252),
    .Y(_13553_));
 sky130_fd_sc_hd__nand3_2 _23506_ (.A(_13548_),
    .B(_06314_),
    .C(_13533_),
    .Y(_13554_));
 sky130_fd_sc_hd__a2bb2oi_4 _23507_ (.A1_N(net284),
    .A2_N(net282),
    .B1(_13533_),
    .B2(_13548_),
    .Y(_13555_));
 sky130_fd_sc_hd__o221ai_4 _23508_ (.A1(net284),
    .A2(net282),
    .B1(_13531_),
    .B2(net240),
    .C1(_13549_),
    .Y(_13556_));
 sky130_fd_sc_hd__nor2_1 _23509_ (.A(_13553_),
    .B(_13555_),
    .Y(_13557_));
 sky130_fd_sc_hd__o211ai_1 _23510_ (.A1(_13128_),
    .A2(_13551_),
    .B1(_13554_),
    .C1(_13556_),
    .Y(_13559_));
 sky130_fd_sc_hd__o2bb2ai_1 _23511_ (.A1_N(_13127_),
    .A2_N(_13138_),
    .B1(_13553_),
    .B2(_13555_),
    .Y(_13560_));
 sky130_fd_sc_hd__nand3_2 _23512_ (.A(_13556_),
    .B(_13552_),
    .C(_13554_),
    .Y(_13561_));
 sky130_fd_sc_hd__o22ai_4 _23513_ (.A1(_13128_),
    .A2(_13551_),
    .B1(_13553_),
    .B2(_13555_),
    .Y(_13562_));
 sky130_fd_sc_hd__nand3_2 _23514_ (.A(_13560_),
    .B(net213),
    .C(_13559_),
    .Y(_13563_));
 sky130_fd_sc_hd__o221a_1 _23515_ (.A1(_06286_),
    .A2(_06288_),
    .B1(_13531_),
    .B2(net240),
    .C1(_13549_),
    .X(_13564_));
 sky130_fd_sc_hd__o211ai_2 _23516_ (.A1(net239),
    .A2(_06292_),
    .B1(_13561_),
    .C1(_13562_),
    .Y(_13565_));
 sky130_fd_sc_hd__o21ai_2 _23517_ (.A1(net213),
    .A2(_13550_),
    .B1(_13563_),
    .Y(_13566_));
 sky130_fd_sc_hd__a311oi_4 _23518_ (.A1(_13561_),
    .A2(_13562_),
    .A3(net213),
    .B1(_13564_),
    .C1(_06014_),
    .Y(_13567_));
 sky130_fd_sc_hd__nand3b_4 _23519_ (.A_N(_13564_),
    .B(_13565_),
    .C(net254),
    .Y(_13568_));
 sky130_fd_sc_hd__o211a_1 _23520_ (.A1(_13550_),
    .A2(net213),
    .B1(_06014_),
    .C1(_13563_),
    .X(_13570_));
 sky130_fd_sc_hd__o211ai_4 _23521_ (.A1(_13550_),
    .A2(net213),
    .B1(_06014_),
    .C1(_13563_),
    .Y(_13571_));
 sky130_fd_sc_hd__nand2_1 _23522_ (.A(_13568_),
    .B(_13571_),
    .Y(_13572_));
 sky130_fd_sc_hd__o2bb2ai_1 _23523_ (.A1_N(_13149_),
    .A2_N(_13150_),
    .B1(net263),
    .B2(_13142_),
    .Y(_13573_));
 sky130_fd_sc_hd__o2bb2ai_1 _23524_ (.A1_N(_13143_),
    .A2_N(_13158_),
    .B1(_13567_),
    .B2(_13570_),
    .Y(_13574_));
 sky130_fd_sc_hd__o2111ai_4 _23525_ (.A1(_13142_),
    .A2(net263),
    .B1(_13568_),
    .C1(_13158_),
    .D1(_13571_),
    .Y(_13575_));
 sky130_fd_sc_hd__o211ai_2 _23526_ (.A1(net263),
    .A2(_13142_),
    .B1(_13158_),
    .C1(_13572_),
    .Y(_13576_));
 sky130_fd_sc_hd__o2111ai_4 _23527_ (.A1(_05768_),
    .A2(_13140_),
    .B1(_13568_),
    .C1(_13571_),
    .D1(_13573_),
    .Y(_13577_));
 sky130_fd_sc_hd__a22oi_4 _23528_ (.A1(_06609_),
    .A2(_06611_),
    .B1(_13574_),
    .B2(_13575_),
    .Y(_13578_));
 sky130_fd_sc_hd__nand3_2 _23529_ (.A(_13576_),
    .B(_13577_),
    .C(net210),
    .Y(_13579_));
 sky130_fd_sc_hd__o211a_1 _23530_ (.A1(_13550_),
    .A2(net213),
    .B1(_06613_),
    .C1(_13563_),
    .X(_13581_));
 sky130_fd_sc_hd__or3_1 _23531_ (.A(net238),
    .B(_06610_),
    .C(_13566_),
    .X(_13582_));
 sky130_fd_sc_hd__o31a_1 _23532_ (.A1(net238),
    .A2(_06610_),
    .A3(_13566_),
    .B1(_13579_),
    .X(_13583_));
 sky130_fd_sc_hd__a31o_1 _23533_ (.A1(_13576_),
    .A2(_13577_),
    .A3(net210),
    .B1(_13581_),
    .X(_13584_));
 sky130_fd_sc_hd__a22oi_1 _23534_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_13579_),
    .B2(_13582_),
    .Y(_13585_));
 sky130_fd_sc_hd__o22ai_4 _23535_ (.A1(_05760_),
    .A2(_05762_),
    .B1(_13578_),
    .B2(_13581_),
    .Y(_13586_));
 sky130_fd_sc_hd__a31oi_1 _23536_ (.A1(_13576_),
    .A2(_13577_),
    .A3(net210),
    .B1(_05768_),
    .Y(_13587_));
 sky130_fd_sc_hd__o221ai_4 _23537_ (.A1(_05765_),
    .A2(_05766_),
    .B1(net210),
    .B2(_13566_),
    .C1(_13579_),
    .Y(_13588_));
 sky130_fd_sc_hd__a21oi_1 _23538_ (.A1(_13582_),
    .A2(_13587_),
    .B1(_13585_),
    .Y(_13589_));
 sky130_fd_sc_hd__nand2_1 _23539_ (.A(_13586_),
    .B(_13588_),
    .Y(_13590_));
 sky130_fd_sc_hd__nand3_1 _23540_ (.A(_12259_),
    .B(_12261_),
    .C(_11795_),
    .Y(_13592_));
 sky130_fd_sc_hd__o21bai_1 _23541_ (.A1(net295),
    .A2(_12686_),
    .B1_N(_13592_),
    .Y(_13593_));
 sky130_fd_sc_hd__nor3_2 _23542_ (.A(_12694_),
    .B(_13592_),
    .C(_12695_),
    .Y(_13594_));
 sky130_fd_sc_hd__nand2_1 _23543_ (.A(_13165_),
    .B(_13594_),
    .Y(_13595_));
 sky130_fd_sc_hd__o211a_1 _23544_ (.A1(_13170_),
    .A2(_13164_),
    .B1(_13166_),
    .C1(_13595_),
    .X(_13596_));
 sky130_fd_sc_hd__o211ai_4 _23545_ (.A1(_13170_),
    .A2(_13164_),
    .B1(_13166_),
    .C1(_13595_),
    .Y(_13597_));
 sky130_fd_sc_hd__nor3_1 _23546_ (.A(_11797_),
    .B(_12694_),
    .C(_13593_),
    .Y(_13598_));
 sky130_fd_sc_hd__o211ai_4 _23547_ (.A1(_11312_),
    .A2(_11796_),
    .B1(_13594_),
    .C1(_13166_),
    .Y(_13599_));
 sky130_fd_sc_hd__nand3_1 _23548_ (.A(_13598_),
    .B(_13166_),
    .C(_13165_),
    .Y(_13600_));
 sky130_fd_sc_hd__o21ai_2 _23549_ (.A1(_13164_),
    .A2(_13599_),
    .B1(_13597_),
    .Y(_13601_));
 sky130_fd_sc_hd__a21oi_1 _23550_ (.A1(_13597_),
    .A2(_13600_),
    .B1(_13590_),
    .Y(_13603_));
 sky130_fd_sc_hd__o22ai_2 _23551_ (.A1(_06899_),
    .A2(net228),
    .B1(_13589_),
    .B2(_13601_),
    .Y(_13604_));
 sky130_fd_sc_hd__and3_1 _23552_ (.A(_06900_),
    .B(_06902_),
    .C(_13584_),
    .X(_13605_));
 sky130_fd_sc_hd__inv_2 _23553_ (.A(_13605_),
    .Y(_13606_));
 sky130_fd_sc_hd__a22o_1 _23554_ (.A1(_13586_),
    .A2(_13588_),
    .B1(_13597_),
    .B2(_13600_),
    .X(_13607_));
 sky130_fd_sc_hd__o31ai_2 _23555_ (.A1(_13581_),
    .A2(_05768_),
    .A3(_13578_),
    .B1(_13600_),
    .Y(_13608_));
 sky130_fd_sc_hd__o211ai_4 _23556_ (.A1(_13599_),
    .A2(_13164_),
    .B1(_13588_),
    .C1(_13597_),
    .Y(_13609_));
 sky130_fd_sc_hd__o2111ai_4 _23557_ (.A1(_13599_),
    .A2(_13164_),
    .B1(_13588_),
    .C1(_13597_),
    .D1(_13586_),
    .Y(_13610_));
 sky130_fd_sc_hd__nand3_2 _23558_ (.A(_13607_),
    .B(_13610_),
    .C(net208),
    .Y(_13611_));
 sky130_fd_sc_hd__a31o_2 _23559_ (.A1(_13607_),
    .A2(_13610_),
    .A3(net208),
    .B1(_13605_),
    .X(_13612_));
 sky130_fd_sc_hd__inv_2 _23560_ (.A(_13612_),
    .Y(_13614_));
 sky130_fd_sc_hd__a211o_2 _23561_ (.A1(_13606_),
    .A2(_13611_),
    .B1(_07227_),
    .C1(net206),
    .X(_13615_));
 sky130_fd_sc_hd__a311oi_2 _23562_ (.A1(_13607_),
    .A2(_13610_),
    .A3(net208),
    .B1(_13605_),
    .C1(net292),
    .Y(_13616_));
 sky130_fd_sc_hd__nand3_4 _23563_ (.A(_13611_),
    .B(_05507_),
    .C(_13606_),
    .Y(_13617_));
 sky130_fd_sc_hd__o221ai_4 _23564_ (.A1(net208),
    .A2(_13584_),
    .B1(_13603_),
    .B2(_13604_),
    .C1(net292),
    .Y(_13618_));
 sky130_fd_sc_hd__o221a_1 _23565_ (.A1(_12708_),
    .A2(_12712_),
    .B1(_13179_),
    .B2(net295),
    .C1(_12707_),
    .X(_13619_));
 sky130_fd_sc_hd__a31o_1 _23566_ (.A1(net294),
    .A2(_13177_),
    .A3(_13178_),
    .B1(_13183_),
    .X(_13620_));
 sky130_fd_sc_hd__o31ai_2 _23567_ (.A1(_12708_),
    .A2(_13182_),
    .A3(_13186_),
    .B1(_13189_),
    .Y(_13621_));
 sky130_fd_sc_hd__a21oi_1 _23568_ (.A1(_13187_),
    .A2(_13183_),
    .B1(_13188_),
    .Y(_13622_));
 sky130_fd_sc_hd__a21oi_1 _23569_ (.A1(_13617_),
    .A2(_13618_),
    .B1(_13621_),
    .Y(_13623_));
 sky130_fd_sc_hd__o2bb2ai_4 _23570_ (.A1_N(_13617_),
    .A2_N(_13618_),
    .B1(_13619_),
    .B2(_13186_),
    .Y(_13625_));
 sky130_fd_sc_hd__o2111a_1 _23571_ (.A1(net294),
    .A2(_13180_),
    .B1(_13617_),
    .C1(_13618_),
    .D1(_13620_),
    .X(_13626_));
 sky130_fd_sc_hd__o2111ai_1 _23572_ (.A1(net294),
    .A2(_13180_),
    .B1(_13617_),
    .C1(_13618_),
    .D1(_13620_),
    .Y(_13627_));
 sky130_fd_sc_hd__a31oi_4 _23573_ (.A1(_13617_),
    .A2(_13618_),
    .A3(_13621_),
    .B1(_07232_),
    .Y(_13628_));
 sky130_fd_sc_hd__nand3_2 _23574_ (.A(net185),
    .B(_13625_),
    .C(_13627_),
    .Y(_13629_));
 sky130_fd_sc_hd__o22ai_2 _23575_ (.A1(_07227_),
    .A2(net206),
    .B1(_13623_),
    .B2(_13626_),
    .Y(_13630_));
 sky130_fd_sc_hd__o31a_1 _23576_ (.A1(_07227_),
    .A2(net206),
    .A3(_13614_),
    .B1(_13629_),
    .X(_13631_));
 sky130_fd_sc_hd__a22o_1 _23577_ (.A1(_07232_),
    .A2(_13612_),
    .B1(_13628_),
    .B2(_13625_),
    .X(_13632_));
 sky130_fd_sc_hd__o211a_1 _23578_ (.A1(_12722_),
    .A2(_12730_),
    .B1(_13201_),
    .C1(_12721_),
    .X(_13633_));
 sky130_fd_sc_hd__o221a_1 _23579_ (.A1(_02148_),
    .A2(_12718_),
    .B1(_04238_),
    .B2(_13198_),
    .C1(_13205_),
    .X(_13634_));
 sky130_fd_sc_hd__o21ai_1 _23580_ (.A1(_13202_),
    .A2(_13206_),
    .B1(_13201_),
    .Y(_13636_));
 sky130_fd_sc_hd__a21oi_1 _23581_ (.A1(_13628_),
    .A2(_13625_),
    .B1(net294),
    .Y(_13637_));
 sky130_fd_sc_hd__a221oi_4 _23582_ (.A1(_07232_),
    .A2(_13612_),
    .B1(_13628_),
    .B2(_13625_),
    .C1(net294),
    .Y(_13638_));
 sky130_fd_sc_hd__o211ai_4 _23583_ (.A1(net185),
    .A2(_13614_),
    .B1(net295),
    .C1(_13629_),
    .Y(_13639_));
 sky130_fd_sc_hd__a2bb2oi_4 _23584_ (.A1_N(net318),
    .A2_N(net316),
    .B1(_13615_),
    .B2(_13629_),
    .Y(_13640_));
 sky130_fd_sc_hd__o221ai_4 _23585_ (.A1(net318),
    .A2(net316),
    .B1(net185),
    .B2(_13612_),
    .C1(_13630_),
    .Y(_13641_));
 sky130_fd_sc_hd__o211ai_2 _23586_ (.A1(_13202_),
    .A2(_13633_),
    .B1(_13639_),
    .C1(_13641_),
    .Y(_13642_));
 sky130_fd_sc_hd__o22ai_2 _23587_ (.A1(_13200_),
    .A2(_13634_),
    .B1(_13638_),
    .B2(_13640_),
    .Y(_13643_));
 sky130_fd_sc_hd__o211ai_4 _23588_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_13642_),
    .C1(_13643_),
    .Y(_13644_));
 sky130_fd_sc_hd__o311a_1 _23589_ (.A1(_07227_),
    .A2(net206),
    .A3(_13612_),
    .B1(_13630_),
    .C1(_07550_),
    .X(_13645_));
 sky130_fd_sc_hd__o211ai_4 _23590_ (.A1(_13200_),
    .A2(_13634_),
    .B1(_13639_),
    .C1(_13641_),
    .Y(_13647_));
 sky130_fd_sc_hd__o22ai_4 _23591_ (.A1(_13202_),
    .A2(_13633_),
    .B1(_13638_),
    .B2(_13640_),
    .Y(_13648_));
 sky130_fd_sc_hd__o211ai_2 _23592_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_13647_),
    .C1(_13648_),
    .Y(_13649_));
 sky130_fd_sc_hd__a31oi_4 _23593_ (.A1(_13648_),
    .A2(net163),
    .A3(_13647_),
    .B1(_13645_),
    .Y(_13650_));
 sky130_fd_sc_hd__o211a_1 _23594_ (.A1(_13632_),
    .A2(net163),
    .B1(_04238_),
    .C1(_13644_),
    .X(_13651_));
 sky130_fd_sc_hd__o211ai_4 _23595_ (.A1(_13632_),
    .A2(net163),
    .B1(_04238_),
    .C1(_13644_),
    .Y(_13652_));
 sky130_fd_sc_hd__o211a_1 _23596_ (.A1(net163),
    .A2(_13631_),
    .B1(_04227_),
    .C1(_13649_),
    .X(_13653_));
 sky130_fd_sc_hd__o211ai_4 _23597_ (.A1(net163),
    .A2(_13631_),
    .B1(_04227_),
    .C1(_13649_),
    .Y(_13654_));
 sky130_fd_sc_hd__o22a_1 _23598_ (.A1(_02137_),
    .A2(_13215_),
    .B1(_13222_),
    .B2(_12742_),
    .X(_13655_));
 sky130_fd_sc_hd__a31o_1 _23599_ (.A1(_12743_),
    .A2(_13221_),
    .A3(_13223_),
    .B1(_13217_),
    .X(_13656_));
 sky130_fd_sc_hd__o2bb2ai_2 _23600_ (.A1_N(_13652_),
    .A2_N(_13654_),
    .B1(_13655_),
    .B2(_13220_),
    .Y(_13658_));
 sky130_fd_sc_hd__nand3_2 _23601_ (.A(_13652_),
    .B(_13654_),
    .C(_13656_),
    .Y(_13659_));
 sky130_fd_sc_hd__nand3_1 _23602_ (.A(_13658_),
    .B(_13659_),
    .C(net161),
    .Y(_13660_));
 sky130_fd_sc_hd__o211a_1 _23603_ (.A1(_13632_),
    .A2(net163),
    .B1(_07917_),
    .C1(_13644_),
    .X(_13661_));
 sky130_fd_sc_hd__or3_1 _23604_ (.A(_07912_),
    .B(_07914_),
    .C(_13650_),
    .X(_13662_));
 sky130_fd_sc_hd__a31o_1 _23605_ (.A1(_13658_),
    .A2(_13659_),
    .A3(net161),
    .B1(_13661_),
    .X(_13663_));
 sky130_fd_sc_hd__a21oi_2 _23606_ (.A1(_13660_),
    .A2(_13662_),
    .B1(_02137_),
    .Y(_13664_));
 sky130_fd_sc_hd__a22o_1 _23607_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_13660_),
    .B2(_13662_),
    .X(_13665_));
 sky130_fd_sc_hd__a311oi_4 _23608_ (.A1(_13658_),
    .A2(_13659_),
    .A3(net161),
    .B1(_13661_),
    .C1(_02148_),
    .Y(_13666_));
 sky130_fd_sc_hd__a311o_2 _23609_ (.A1(_13658_),
    .A2(_13659_),
    .A3(net161),
    .B1(_13661_),
    .C1(_02148_),
    .X(_13667_));
 sky130_fd_sc_hd__nand4_2 _23610_ (.A(_11860_),
    .B(_11862_),
    .C(_12324_),
    .D(_12326_),
    .Y(_13669_));
 sky130_fd_sc_hd__a21oi_2 _23611_ (.A1(_12899_),
    .A2(_12756_),
    .B1(_13669_),
    .Y(_13670_));
 sky130_fd_sc_hd__a211oi_2 _23612_ (.A1(_12761_),
    .A2(_12740_),
    .B1(_13669_),
    .C1(_12764_),
    .Y(_13671_));
 sky130_fd_sc_hd__nand3_1 _23613_ (.A(_13670_),
    .B(_13238_),
    .C(_12763_),
    .Y(_13672_));
 sky130_fd_sc_hd__nand4_1 _23614_ (.A(_12763_),
    .B(_13670_),
    .C(_13238_),
    .D(_11864_),
    .Y(_13673_));
 sky130_fd_sc_hd__o221ai_4 _23615_ (.A1(_13234_),
    .A2(_00251_),
    .B1(_13671_),
    .B2(_13247_),
    .C1(_13673_),
    .Y(_13674_));
 sky130_fd_sc_hd__o211ai_4 _23616_ (.A1(_13237_),
    .A2(_13245_),
    .B1(_13672_),
    .C1(_13241_),
    .Y(_13675_));
 sky130_fd_sc_hd__o2111ai_4 _23617_ (.A1(_12899_),
    .A2(_12756_),
    .B1(_13238_),
    .C1(_13670_),
    .D1(_13241_),
    .Y(_13676_));
 sky130_fd_sc_hd__nand4_2 _23618_ (.A(_13238_),
    .B(_13671_),
    .C(_13241_),
    .D(_11864_),
    .Y(_13677_));
 sky130_fd_sc_hd__o21ai_2 _23619_ (.A1(_11865_),
    .A2(_13676_),
    .B1(_13675_),
    .Y(_13678_));
 sky130_fd_sc_hd__inv_2 _23620_ (.A(_13678_),
    .Y(_13680_));
 sky130_fd_sc_hd__o221ai_2 _23621_ (.A1(_13233_),
    .A2(_00240_),
    .B1(_13666_),
    .B2(_13664_),
    .C1(_13674_),
    .Y(_13681_));
 sky130_fd_sc_hd__nand4_1 _23622_ (.A(_13665_),
    .B(_13667_),
    .C(_13675_),
    .D(_13677_),
    .Y(_13682_));
 sky130_fd_sc_hd__o2111ai_1 _23623_ (.A1(_00240_),
    .A2(_13233_),
    .B1(_13665_),
    .C1(_13667_),
    .D1(_13674_),
    .Y(_13683_));
 sky130_fd_sc_hd__o221ai_2 _23624_ (.A1(_11865_),
    .A2(_13676_),
    .B1(_13666_),
    .B2(_13664_),
    .C1(_13675_),
    .Y(_13684_));
 sky130_fd_sc_hd__nand3_2 _23625_ (.A(_13683_),
    .B(_13684_),
    .C(_08300_),
    .Y(_13685_));
 sky130_fd_sc_hd__and3_1 _23626_ (.A(_08297_),
    .B(_08299_),
    .C(_13663_),
    .X(_13686_));
 sky130_fd_sc_hd__a211o_1 _23627_ (.A1(_13660_),
    .A2(_13662_),
    .B1(net180),
    .C1(_08298_),
    .X(_13687_));
 sky130_fd_sc_hd__nand3_2 _23628_ (.A(_13681_),
    .B(_13682_),
    .C(_08300_),
    .Y(_13688_));
 sky130_fd_sc_hd__o311a_2 _23629_ (.A1(net180),
    .A2(_13663_),
    .A3(_08298_),
    .B1(_08715_),
    .C1(_13685_),
    .X(_13689_));
 sky130_fd_sc_hd__a22o_2 _23630_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_13687_),
    .B2(_13688_),
    .X(_13691_));
 sky130_fd_sc_hd__a31o_1 _23631_ (.A1(_13681_),
    .A2(_13682_),
    .A3(_08300_),
    .B1(_00251_),
    .X(_13692_));
 sky130_fd_sc_hd__o211ai_4 _23632_ (.A1(_00218_),
    .A2(_00229_),
    .B1(_13687_),
    .C1(_13688_),
    .Y(_13693_));
 sky130_fd_sc_hd__a2bb2oi_1 _23633_ (.A1_N(_00174_),
    .A2_N(net344),
    .B1(_13687_),
    .B2(_13688_),
    .Y(_13694_));
 sky130_fd_sc_hd__o211ai_4 _23634_ (.A1(_13663_),
    .A2(_08300_),
    .B1(_00251_),
    .C1(_13685_),
    .Y(_13695_));
 sky130_fd_sc_hd__o211a_1 _23635_ (.A1(_12781_),
    .A2(_12784_),
    .B1(_13260_),
    .C1(_12780_),
    .X(_13696_));
 sky130_fd_sc_hd__o32a_2 _23636_ (.A1(net361),
    .A2(net345),
    .A3(_13252_),
    .B1(_13256_),
    .B2(_13259_),
    .X(_13697_));
 sky130_fd_sc_hd__o2bb2ai_4 _23637_ (.A1_N(_13693_),
    .A2_N(_13695_),
    .B1(_13696_),
    .B2(_13257_),
    .Y(_13698_));
 sky130_fd_sc_hd__nand3_4 _23638_ (.A(_13693_),
    .B(_13695_),
    .C(_13697_),
    .Y(_13699_));
 sky130_fd_sc_hd__nand3_2 _23639_ (.A(_13698_),
    .B(_13699_),
    .C(_08714_),
    .Y(_13700_));
 sky130_fd_sc_hd__a31oi_4 _23640_ (.A1(_13698_),
    .A2(_13699_),
    .A3(_08714_),
    .B1(_13689_),
    .Y(_13702_));
 sky130_fd_sc_hd__a311o_1 _23641_ (.A1(_13698_),
    .A2(_13699_),
    .A3(_08714_),
    .B1(_09125_),
    .C1(_13689_),
    .X(_13703_));
 sky130_fd_sc_hd__o21ai_2 _23642_ (.A1(_12794_),
    .A2(_13275_),
    .B1(_13271_),
    .Y(_13704_));
 sky130_fd_sc_hd__o21ai_2 _23643_ (.A1(_13276_),
    .A2(_13272_),
    .B1(_13271_),
    .Y(_13705_));
 sky130_fd_sc_hd__a31o_1 _23644_ (.A1(_12793_),
    .A2(_12802_),
    .A3(_13271_),
    .B1(_13272_),
    .X(_13706_));
 sky130_fd_sc_hd__a311oi_4 _23645_ (.A1(_13698_),
    .A2(_13699_),
    .A3(_08714_),
    .B1(_13689_),
    .C1(_12899_),
    .Y(_13707_));
 sky130_fd_sc_hd__o211ai_4 _23646_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_13691_),
    .C1(_13700_),
    .Y(_13708_));
 sky130_fd_sc_hd__a2bb2oi_4 _23647_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_13691_),
    .B2(_13700_),
    .Y(_13709_));
 sky130_fd_sc_hd__a2bb2o_1 _23648_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_13691_),
    .B2(_13700_),
    .X(_13710_));
 sky130_fd_sc_hd__nor2_1 _23649_ (.A(_13707_),
    .B(_13709_),
    .Y(_13711_));
 sky130_fd_sc_hd__nand3_1 _23650_ (.A(_13706_),
    .B(_13708_),
    .C(_13710_),
    .Y(_13713_));
 sky130_fd_sc_hd__o21ai_1 _23651_ (.A1(_13707_),
    .A2(_13709_),
    .B1(_13705_),
    .Y(_13714_));
 sky130_fd_sc_hd__o211ai_2 _23652_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_13713_),
    .C1(_13714_),
    .Y(_13715_));
 sky130_fd_sc_hd__or3_1 _23653_ (.A(_09120_),
    .B(_09121_),
    .C(_13702_),
    .X(_13716_));
 sky130_fd_sc_hd__o21ai_1 _23654_ (.A1(_12888_),
    .A2(_13702_),
    .B1(_13705_),
    .Y(_13717_));
 sky130_fd_sc_hd__o2111ai_1 _23655_ (.A1(_11309_),
    .A2(_13270_),
    .B1(_13704_),
    .C1(_13708_),
    .D1(_13710_),
    .Y(_13718_));
 sky130_fd_sc_hd__o2bb2ai_2 _23656_ (.A1_N(_13274_),
    .A2_N(_13704_),
    .B1(_13707_),
    .B2(_13709_),
    .Y(_13719_));
 sky130_fd_sc_hd__o221ai_4 _23657_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_13707_),
    .B2(_13717_),
    .C1(_13719_),
    .Y(_13720_));
 sky130_fd_sc_hd__o21ai_4 _23658_ (.A1(_09125_),
    .A2(_13702_),
    .B1(_13720_),
    .Y(_13721_));
 sky130_fd_sc_hd__inv_2 _23659_ (.A(_13721_),
    .Y(_13722_));
 sky130_fd_sc_hd__a2bb2oi_1 _23660_ (.A1_N(_11210_),
    .A2_N(_11232_),
    .B1(_13716_),
    .B2(_13720_),
    .Y(_13724_));
 sky130_fd_sc_hd__o211ai_4 _23661_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_13703_),
    .C1(_13715_),
    .Y(_13725_));
 sky130_fd_sc_hd__a31oi_1 _23662_ (.A1(_09125_),
    .A2(_13718_),
    .A3(_13719_),
    .B1(_11309_),
    .Y(_13726_));
 sky130_fd_sc_hd__o211a_1 _23663_ (.A1(_09125_),
    .A2(_13702_),
    .B1(_11298_),
    .C1(_13720_),
    .X(_13727_));
 sky130_fd_sc_hd__o211ai_4 _23664_ (.A1(_09125_),
    .A2(_13702_),
    .B1(_11298_),
    .C1(_13720_),
    .Y(_13728_));
 sky130_fd_sc_hd__nand2_2 _23665_ (.A(_13287_),
    .B(_13296_),
    .Y(_13729_));
 sky130_fd_sc_hd__a32o_1 _23666_ (.A1(_10015_),
    .A2(_13280_),
    .A3(_13283_),
    .B1(_13291_),
    .B2(_13287_),
    .X(_13730_));
 sky130_fd_sc_hd__nand3_1 _23667_ (.A(_13725_),
    .B(_13728_),
    .C(_13730_),
    .Y(_13731_));
 sky130_fd_sc_hd__o2bb2ai_1 _23668_ (.A1_N(_13287_),
    .A2_N(_13296_),
    .B1(_13724_),
    .B2(_13727_),
    .Y(_13732_));
 sky130_fd_sc_hd__o2111ai_4 _23669_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .C1(_13731_),
    .D1(_13732_),
    .Y(_13733_));
 sky130_fd_sc_hd__a211o_1 _23670_ (.A1(_13716_),
    .A2(_13720_),
    .B1(_09553_),
    .C1(net155),
    .X(_13735_));
 sky130_fd_sc_hd__inv_2 _23671_ (.A(_13735_),
    .Y(_13736_));
 sky130_fd_sc_hd__a21oi_4 _23672_ (.A1(_13725_),
    .A2(_13728_),
    .B1(_13729_),
    .Y(_13737_));
 sky130_fd_sc_hd__a31o_2 _23673_ (.A1(_13725_),
    .A2(_13729_),
    .A3(_13728_),
    .B1(_09562_),
    .X(_13738_));
 sky130_fd_sc_hd__o21ai_4 _23674_ (.A1(_13737_),
    .A2(_13738_),
    .B1(_13735_),
    .Y(_13739_));
 sky130_fd_sc_hd__and3_1 _23675_ (.A(_13739_),
    .B(_10004_),
    .C(_09982_),
    .X(_13740_));
 sky130_fd_sc_hd__o2111ai_4 _23676_ (.A1(_13721_),
    .A2(net143),
    .B1(_10004_),
    .C1(_09982_),
    .D1(_13733_),
    .Y(_13741_));
 sky130_fd_sc_hd__o21ai_2 _23677_ (.A1(_13737_),
    .A2(_13738_),
    .B1(_10015_),
    .Y(_13742_));
 sky130_fd_sc_hd__o221ai_4 _23678_ (.A1(net143),
    .A2(_13722_),
    .B1(_13737_),
    .B2(_13738_),
    .C1(_10015_),
    .Y(_13743_));
 sky130_fd_sc_hd__o32a_4 _23679_ (.A1(_08863_),
    .A2(_08885_),
    .A3(_13297_),
    .B1(_13298_),
    .B2(_12879_),
    .X(_13744_));
 sky130_fd_sc_hd__o21ai_1 _23680_ (.A1(_12879_),
    .A2(_13298_),
    .B1(_13301_),
    .Y(_13746_));
 sky130_fd_sc_hd__a21oi_2 _23681_ (.A1(_13741_),
    .A2(_13743_),
    .B1(_13744_),
    .Y(_13747_));
 sky130_fd_sc_hd__a31o_1 _23682_ (.A1(_13741_),
    .A2(_13744_),
    .A3(_13743_),
    .B1(_09578_),
    .X(_13748_));
 sky130_fd_sc_hd__or3b_1 _23683_ (.A(_09571_),
    .B(_09573_),
    .C_N(_13739_),
    .X(_13749_));
 sky130_fd_sc_hd__a21o_1 _23684_ (.A1(_13741_),
    .A2(_13743_),
    .B1(_13746_),
    .X(_13750_));
 sky130_fd_sc_hd__o21ai_2 _23685_ (.A1(_10025_),
    .A2(_13739_),
    .B1(_13746_),
    .Y(_13751_));
 sky130_fd_sc_hd__o221ai_4 _23686_ (.A1(_09571_),
    .A2(_09573_),
    .B1(_13740_),
    .B2(_13751_),
    .C1(_13750_),
    .Y(_13752_));
 sky130_fd_sc_hd__o22a_1 _23687_ (.A1(_09579_),
    .A2(_13739_),
    .B1(_13747_),
    .B2(_13748_),
    .X(_13753_));
 sky130_fd_sc_hd__a31oi_2 _23688_ (.A1(_12840_),
    .A2(_13309_),
    .A3(_13310_),
    .B1(_13307_),
    .Y(_13754_));
 sky130_fd_sc_hd__a31o_1 _23689_ (.A1(_12840_),
    .A2(_13309_),
    .A3(_13310_),
    .B1(_13307_),
    .X(_13755_));
 sky130_fd_sc_hd__o211ai_2 _23690_ (.A1(_08863_),
    .A2(_08885_),
    .B1(_13749_),
    .C1(_13752_),
    .Y(_13757_));
 sky130_fd_sc_hd__o221ai_4 _23691_ (.A1(_09579_),
    .A2(_13739_),
    .B1(_13747_),
    .B2(_13748_),
    .C1(_08918_),
    .Y(_13758_));
 sky130_fd_sc_hd__a21oi_1 _23692_ (.A1(_13757_),
    .A2(_13758_),
    .B1(_13754_),
    .Y(_13759_));
 sky130_fd_sc_hd__a31o_1 _23693_ (.A1(_13757_),
    .A2(_13758_),
    .A3(_13754_),
    .B1(_10479_),
    .X(_13760_));
 sky130_fd_sc_hd__o22ai_4 _23694_ (.A1(_10480_),
    .A2(_13753_),
    .B1(_13759_),
    .B2(_13760_),
    .Y(_13761_));
 sky130_fd_sc_hd__a21o_1 _23695_ (.A1(_07811_),
    .A2(_07833_),
    .B1(_13761_),
    .X(_13762_));
 sky130_fd_sc_hd__inv_2 _23696_ (.A(_13762_),
    .Y(_13763_));
 sky130_fd_sc_hd__o21ai_2 _23697_ (.A1(net368),
    .A2(_07866_),
    .B1(_13761_),
    .Y(_13764_));
 sky130_fd_sc_hd__a311o_1 _23698_ (.A1(_13316_),
    .A2(_07022_),
    .A3(net376),
    .B1(_12850_),
    .C1(_12857_),
    .X(_13765_));
 sky130_fd_sc_hd__or3_1 _23699_ (.A(_10949_),
    .B(net136),
    .C(_13761_),
    .X(_13766_));
 sky130_fd_sc_hd__a22o_1 _23700_ (.A1(_13762_),
    .A2(_13764_),
    .B1(_13765_),
    .B2(_13318_),
    .X(_13768_));
 sky130_fd_sc_hd__o211ai_4 _23701_ (.A1(_07044_),
    .A2(_13316_),
    .B1(_13764_),
    .C1(_13765_),
    .Y(_13769_));
 sky130_fd_sc_hd__o221ai_4 _23702_ (.A1(_10949_),
    .A2(net136),
    .B1(_13769_),
    .B2(_13763_),
    .C1(_13768_),
    .Y(_13770_));
 sky130_fd_sc_hd__o21ai_1 _23703_ (.A1(_10954_),
    .A2(_13761_),
    .B1(_13770_),
    .Y(_13771_));
 sky130_fd_sc_hd__o21ai_1 _23704_ (.A1(_06332_),
    .A2(_13324_),
    .B1(_13331_),
    .Y(_13772_));
 sky130_fd_sc_hd__o221ai_4 _23705_ (.A1(_06989_),
    .A2(net375),
    .B1(_10954_),
    .B2(_13761_),
    .C1(_13770_),
    .Y(_13773_));
 sky130_fd_sc_hd__a21oi_1 _23706_ (.A1(_13766_),
    .A2(_13770_),
    .B1(_07033_),
    .Y(_13774_));
 sky130_fd_sc_hd__a22o_1 _23707_ (.A1(_06956_),
    .A2(_06978_),
    .B1(_13766_),
    .B2(_13770_),
    .X(_13775_));
 sky130_fd_sc_hd__a22oi_1 _23708_ (.A1(_13325_),
    .A2(_13331_),
    .B1(_13773_),
    .B2(_13775_),
    .Y(_13776_));
 sky130_fd_sc_hd__a41o_1 _23709_ (.A1(_13325_),
    .A2(_13331_),
    .A3(_13773_),
    .A4(_13775_),
    .B1(_11464_),
    .X(_13777_));
 sky130_fd_sc_hd__o22a_1 _23710_ (.A1(_11465_),
    .A2(_13771_),
    .B1(_13776_),
    .B2(_13777_),
    .X(_13779_));
 sky130_fd_sc_hd__a21oi_1 _23711_ (.A1(_06300_),
    .A2(_06321_),
    .B1(_13779_),
    .Y(_13780_));
 sky130_fd_sc_hd__o221a_1 _23712_ (.A1(_11465_),
    .A2(_13771_),
    .B1(_13776_),
    .B2(_13777_),
    .C1(_06343_),
    .X(_13781_));
 sky130_fd_sc_hd__nor2_1 _23713_ (.A(_13780_),
    .B(_13781_),
    .Y(_13782_));
 sky130_fd_sc_hd__a21o_1 _23714_ (.A1(_13334_),
    .A2(_13336_),
    .B1(_13337_),
    .X(_13783_));
 sky130_fd_sc_hd__o21a_1 _23715_ (.A1(_13783_),
    .A2(_13782_),
    .B1(_11943_),
    .X(_13784_));
 sky130_fd_sc_hd__or2_1 _23716_ (.A(_13779_),
    .B(_13784_),
    .X(_13785_));
 sky130_fd_sc_hd__a21oi_1 _23717_ (.A1(_05119_),
    .A2(_13340_),
    .B1(_13785_),
    .Y(_13786_));
 sky130_fd_sc_hd__and3_1 _23718_ (.A(_05119_),
    .B(_13340_),
    .C(_13785_),
    .X(_13787_));
 sky130_fd_sc_hd__nor2_1 _23719_ (.A(_13786_),
    .B(_13787_),
    .Y(net93));
 sky130_fd_sc_hd__o21ai_1 _23720_ (.A1(_13340_),
    .A2(_13785_),
    .B1(_05119_),
    .Y(_13789_));
 sky130_fd_sc_hd__o311a_1 _23721_ (.A1(_06848_),
    .A2(_10970_),
    .A3(_13341_),
    .B1(_13348_),
    .C1(_11471_),
    .X(_13790_));
 sky130_fd_sc_hd__o311ai_4 _23722_ (.A1(_06848_),
    .A2(_10970_),
    .A3(_13341_),
    .B1(_13348_),
    .C1(_11471_),
    .Y(_13791_));
 sky130_fd_sc_hd__o21ai_1 _23723_ (.A1(net374),
    .A2(_07702_),
    .B1(_13791_),
    .Y(_13792_));
 sky130_fd_sc_hd__or4_1 _23724_ (.A(_07724_),
    .B(_08678_),
    .C(_08700_),
    .D(_13790_),
    .X(_13793_));
 sky130_fd_sc_hd__o211ai_2 _23725_ (.A1(net374),
    .A2(_07702_),
    .B1(_10971_),
    .C1(_13791_),
    .Y(_13794_));
 sky130_fd_sc_hd__a22o_1 _23726_ (.A1(_10966_),
    .A2(_10968_),
    .B1(_13791_),
    .B2(net355),
    .X(_13795_));
 sky130_fd_sc_hd__and2_1 _23727_ (.A(_13794_),
    .B(_13795_),
    .X(_13796_));
 sky130_fd_sc_hd__nand2_1 _23728_ (.A(_13794_),
    .B(_13795_),
    .Y(_13797_));
 sky130_fd_sc_hd__o21bai_1 _23729_ (.A1(_13358_),
    .A2(_13361_),
    .B1_N(_13355_),
    .Y(_13798_));
 sky130_fd_sc_hd__nand2_2 _23730_ (.A(_13798_),
    .B(_13796_),
    .Y(_13800_));
 sky130_fd_sc_hd__o211ai_2 _23731_ (.A1(_13358_),
    .A2(_13361_),
    .B1(_13797_),
    .C1(_13356_),
    .Y(_13801_));
 sky130_fd_sc_hd__nand3_1 _23732_ (.A(_13800_),
    .B(_13801_),
    .C(net338),
    .Y(_13802_));
 sky130_fd_sc_hd__and3_1 _23733_ (.A(_08689_),
    .B(_08711_),
    .C(_13792_),
    .X(_13803_));
 sky130_fd_sc_hd__a22oi_2 _23734_ (.A1(_08689_),
    .A2(_08711_),
    .B1(_13800_),
    .B2(_13801_),
    .Y(_13804_));
 sky130_fd_sc_hd__a21oi_2 _23735_ (.A1(_13793_),
    .A2(_13802_),
    .B1(net335),
    .Y(_13805_));
 sky130_fd_sc_hd__a2bb2oi_1 _23736_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_13793_),
    .B2(_13802_),
    .Y(_13806_));
 sky130_fd_sc_hd__or3_1 _23737_ (.A(net150),
    .B(_13803_),
    .C(_13804_),
    .X(_13807_));
 sky130_fd_sc_hd__a31oi_1 _23738_ (.A1(_13800_),
    .A2(_13801_),
    .A3(net338),
    .B1(_10492_),
    .Y(_13808_));
 sky130_fd_sc_hd__o311a_1 _23739_ (.A1(_07724_),
    .A2(net338),
    .A3(_13790_),
    .B1(net150),
    .C1(_13802_),
    .X(_13809_));
 sky130_fd_sc_hd__o21ai_1 _23740_ (.A1(net338),
    .A2(_13792_),
    .B1(_13808_),
    .Y(_13811_));
 sky130_fd_sc_hd__a21oi_1 _23741_ (.A1(_13793_),
    .A2(_13808_),
    .B1(_13806_),
    .Y(_13812_));
 sky130_fd_sc_hd__o41ai_2 _23742_ (.A1(_10489_),
    .A2(_10490_),
    .A3(_13803_),
    .A4(_13804_),
    .B1(_13811_),
    .Y(_13813_));
 sky130_fd_sc_hd__a21oi_2 _23743_ (.A1(_13373_),
    .A2(_13379_),
    .B1(_13369_),
    .Y(_13814_));
 sky130_fd_sc_hd__o21ai_1 _23744_ (.A1(_13372_),
    .A2(_13378_),
    .B1(_13370_),
    .Y(_13815_));
 sky130_fd_sc_hd__o221ai_2 _23745_ (.A1(_10026_),
    .A2(_13366_),
    .B1(_13806_),
    .B2(_13809_),
    .C1(_13381_),
    .Y(_13816_));
 sky130_fd_sc_hd__nand2_1 _23746_ (.A(_13815_),
    .B(_13812_),
    .Y(_13817_));
 sky130_fd_sc_hd__o221a_2 _23747_ (.A1(net351),
    .A2(_09807_),
    .B1(_13813_),
    .B2(_13814_),
    .C1(_13816_),
    .X(_13818_));
 sky130_fd_sc_hd__o221ai_2 _23748_ (.A1(net351),
    .A2(_09807_),
    .B1(_13813_),
    .B2(_13814_),
    .C1(_13816_),
    .Y(_13819_));
 sky130_fd_sc_hd__o21a_1 _23749_ (.A1(_13805_),
    .A2(_13818_),
    .B1(_11079_),
    .X(_13820_));
 sky130_fd_sc_hd__o21ai_2 _23750_ (.A1(_13805_),
    .A2(_13818_),
    .B1(_11079_),
    .Y(_13822_));
 sky130_fd_sc_hd__o22a_1 _23751_ (.A1(net170),
    .A2(net169),
    .B1(_13805_),
    .B2(_13818_),
    .X(_13823_));
 sky130_fd_sc_hd__o22ai_2 _23752_ (.A1(net170),
    .A2(net169),
    .B1(_13805_),
    .B2(_13818_),
    .Y(_13824_));
 sky130_fd_sc_hd__nand3b_2 _23753_ (.A_N(_13805_),
    .B(_13819_),
    .C(_10026_),
    .Y(_13825_));
 sky130_fd_sc_hd__nand2_1 _23754_ (.A(_13824_),
    .B(_13825_),
    .Y(_13826_));
 sky130_fd_sc_hd__o211a_1 _23755_ (.A1(net177),
    .A2(_12495_),
    .B1(_12065_),
    .C1(_12062_),
    .X(_13827_));
 sky130_fd_sc_hd__and4_1 _23756_ (.A(_12951_),
    .B(_13827_),
    .C(_12953_),
    .D(_12500_),
    .X(_13828_));
 sky130_fd_sc_hd__nand4_2 _23757_ (.A(_12951_),
    .B(_13827_),
    .C(_12953_),
    .D(_12500_),
    .Y(_13829_));
 sky130_fd_sc_hd__o211ai_4 _23758_ (.A1(_13829_),
    .A2(_13390_),
    .B1(_13389_),
    .C1(_13392_),
    .Y(_13830_));
 sky130_fd_sc_hd__nand4_4 _23759_ (.A(_13389_),
    .B(_13828_),
    .C(_13391_),
    .D(_12060_),
    .Y(_13831_));
 sky130_fd_sc_hd__nand2_1 _23760_ (.A(_13830_),
    .B(_13831_),
    .Y(_13833_));
 sky130_fd_sc_hd__a22o_1 _23761_ (.A1(_13824_),
    .A2(_13825_),
    .B1(_13830_),
    .B2(_13831_),
    .X(_13834_));
 sky130_fd_sc_hd__nand4_2 _23762_ (.A(_13824_),
    .B(_13825_),
    .C(_13830_),
    .D(_13831_),
    .Y(_13835_));
 sky130_fd_sc_hd__o221a_1 _23763_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_13826_),
    .B2(_13833_),
    .C1(_13834_),
    .X(_13836_));
 sky130_fd_sc_hd__nand3_2 _23764_ (.A(_13834_),
    .B(_13835_),
    .C(net332),
    .Y(_13837_));
 sky130_fd_sc_hd__a21oi_2 _23765_ (.A1(_13822_),
    .A2(_13837_),
    .B1(net311),
    .Y(_13838_));
 sky130_fd_sc_hd__a211o_2 _23766_ (.A1(_13822_),
    .A2(_13837_),
    .B1(net329),
    .C1(net327),
    .X(_13839_));
 sky130_fd_sc_hd__a21oi_1 _23767_ (.A1(_12970_),
    .A2(_13402_),
    .B1(_13397_),
    .Y(_13840_));
 sky130_fd_sc_hd__a31o_1 _23768_ (.A1(_12970_),
    .A2(_13400_),
    .A3(_13402_),
    .B1(_13397_),
    .X(_13841_));
 sky130_fd_sc_hd__a31oi_2 _23769_ (.A1(_12970_),
    .A2(_13400_),
    .A3(_13402_),
    .B1(_13397_),
    .Y(_13842_));
 sky130_fd_sc_hd__a311oi_4 _23770_ (.A1(_13834_),
    .A2(_13835_),
    .A3(net332),
    .B1(_09595_),
    .C1(_13820_),
    .Y(_13844_));
 sky130_fd_sc_hd__nand3_2 _23771_ (.A(_13837_),
    .B(net172),
    .C(_13822_),
    .Y(_13845_));
 sky130_fd_sc_hd__a2bb2oi_1 _23772_ (.A1_N(_09588_),
    .A2_N(_09590_),
    .B1(_13822_),
    .B2(_13837_),
    .Y(_13846_));
 sky130_fd_sc_hd__o22ai_4 _23773_ (.A1(_09588_),
    .A2(_09590_),
    .B1(_13820_),
    .B2(_13836_),
    .Y(_13847_));
 sky130_fd_sc_hd__nand3_4 _23774_ (.A(_13847_),
    .B(_13841_),
    .C(_13845_),
    .Y(_13848_));
 sky130_fd_sc_hd__o22ai_4 _23775_ (.A1(_13399_),
    .A2(_13840_),
    .B1(_13844_),
    .B2(_13846_),
    .Y(_13849_));
 sky130_fd_sc_hd__o211ai_4 _23776_ (.A1(net329),
    .A2(net327),
    .B1(_13848_),
    .C1(_13849_),
    .Y(_13850_));
 sky130_fd_sc_hd__a31o_1 _23777_ (.A1(_13848_),
    .A2(_13849_),
    .A3(net311),
    .B1(_13838_),
    .X(_13851_));
 sky130_fd_sc_hd__o211ai_4 _23778_ (.A1(net199),
    .A2(_12978_),
    .B1(_13413_),
    .C1(_13417_),
    .Y(_13852_));
 sky130_fd_sc_hd__o21ai_1 _23779_ (.A1(net175),
    .A2(_13412_),
    .B1(_13852_),
    .Y(_13853_));
 sky130_fd_sc_hd__a311oi_4 _23780_ (.A1(_13848_),
    .A2(_13849_),
    .A3(net311),
    .B1(net173),
    .C1(_13838_),
    .Y(_13855_));
 sky130_fd_sc_hd__nand3_2 _23781_ (.A(_13850_),
    .B(net174),
    .C(_13839_),
    .Y(_13856_));
 sky130_fd_sc_hd__a2bb2oi_4 _23782_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_13839_),
    .B2(_13850_),
    .Y(_13857_));
 sky130_fd_sc_hd__a2bb2o_1 _23783_ (.A1_N(_09134_),
    .A2_N(net193),
    .B1(_13839_),
    .B2(_13850_),
    .X(_13858_));
 sky130_fd_sc_hd__nor2_1 _23784_ (.A(_13855_),
    .B(_13857_),
    .Y(_13859_));
 sky130_fd_sc_hd__nand3_1 _23785_ (.A(_13853_),
    .B(_13856_),
    .C(_13858_),
    .Y(_13860_));
 sky130_fd_sc_hd__o221ai_4 _23786_ (.A1(net175),
    .A2(_13412_),
    .B1(_13855_),
    .B2(_13857_),
    .C1(_13852_),
    .Y(_13861_));
 sky130_fd_sc_hd__o211ai_4 _23787_ (.A1(_00011_),
    .A2(net321),
    .B1(_13860_),
    .C1(_13861_),
    .Y(_13862_));
 sky130_fd_sc_hd__a211o_2 _23788_ (.A1(_13839_),
    .A2(_13850_),
    .B1(_00011_),
    .C1(net321),
    .X(_13863_));
 sky130_fd_sc_hd__o2111ai_4 _23789_ (.A1(net175),
    .A2(_13412_),
    .B1(_13852_),
    .C1(_13856_),
    .D1(_13858_),
    .Y(_13864_));
 sky130_fd_sc_hd__o21ai_1 _23790_ (.A1(_13855_),
    .A2(_13857_),
    .B1(_13853_),
    .Y(_13866_));
 sky130_fd_sc_hd__o211ai_4 _23791_ (.A1(_00011_),
    .A2(net321),
    .B1(_13864_),
    .C1(_13866_),
    .Y(_13867_));
 sky130_fd_sc_hd__o21a_2 _23792_ (.A1(net307),
    .A2(_13851_),
    .B1(_13862_),
    .X(_13868_));
 sky130_fd_sc_hd__and3_2 _23793_ (.A(_01973_),
    .B(_13863_),
    .C(_13867_),
    .X(_13869_));
 sky130_fd_sc_hd__o211ai_4 _23794_ (.A1(_13851_),
    .A2(net307),
    .B1(net175),
    .C1(_13862_),
    .Y(_13870_));
 sky130_fd_sc_hd__o211ai_4 _23795_ (.A1(_08728_),
    .A2(net195),
    .B1(_13863_),
    .C1(_13867_),
    .Y(_13871_));
 sky130_fd_sc_hd__nand2_1 _23796_ (.A(_13870_),
    .B(_13871_),
    .Y(_13872_));
 sky130_fd_sc_hd__a22o_1 _23797_ (.A1(net198),
    .A2(_13424_),
    .B1(_13439_),
    .B2(_13441_),
    .X(_13873_));
 sky130_fd_sc_hd__o211ai_4 _23798_ (.A1(_13430_),
    .A2(_13422_),
    .B1(_13441_),
    .C1(_13439_),
    .Y(_13874_));
 sky130_fd_sc_hd__o2111ai_4 _23799_ (.A1(net199),
    .A2(_13423_),
    .B1(_13870_),
    .C1(_13871_),
    .D1(_13874_),
    .Y(_13875_));
 sky130_fd_sc_hd__o221ai_4 _23800_ (.A1(_13430_),
    .A2(_13422_),
    .B1(_13428_),
    .B2(_13442_),
    .C1(_13872_),
    .Y(_13877_));
 sky130_fd_sc_hd__o211ai_2 _23801_ (.A1(net304),
    .A2(_01951_),
    .B1(_13875_),
    .C1(_13877_),
    .Y(_13878_));
 sky130_fd_sc_hd__a211o_1 _23802_ (.A1(_13863_),
    .A2(_13867_),
    .B1(net304),
    .C1(_01951_),
    .X(_13879_));
 sky130_fd_sc_hd__o2111ai_4 _23803_ (.A1(net198),
    .A2(_13424_),
    .B1(_13870_),
    .C1(_13871_),
    .D1(_13873_),
    .Y(_13880_));
 sky130_fd_sc_hd__o221ai_2 _23804_ (.A1(net199),
    .A2(_13423_),
    .B1(_13433_),
    .B2(_13443_),
    .C1(_13872_),
    .Y(_13881_));
 sky130_fd_sc_hd__nand3_1 _23805_ (.A(_13880_),
    .B(_13881_),
    .C(net278),
    .Y(_13882_));
 sky130_fd_sc_hd__a31oi_4 _23806_ (.A1(_13877_),
    .A2(net278),
    .A3(_13875_),
    .B1(_13869_),
    .Y(_13883_));
 sky130_fd_sc_hd__a31o_1 _23807_ (.A1(_13877_),
    .A2(net278),
    .A3(_13875_),
    .B1(_13869_),
    .X(_13884_));
 sky130_fd_sc_hd__a311oi_4 _23808_ (.A1(_13877_),
    .A2(net278),
    .A3(_13875_),
    .B1(net199),
    .C1(_13869_),
    .Y(_13885_));
 sky130_fd_sc_hd__o211ai_2 _23809_ (.A1(net278),
    .A2(_13868_),
    .B1(_13878_),
    .C1(net198),
    .Y(_13886_));
 sky130_fd_sc_hd__a31oi_1 _23810_ (.A1(_13880_),
    .A2(_13881_),
    .A3(net278),
    .B1(net198),
    .Y(_13888_));
 sky130_fd_sc_hd__o211ai_4 _23811_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_13879_),
    .C1(_13882_),
    .Y(_13889_));
 sky130_fd_sc_hd__a21oi_2 _23812_ (.A1(_13888_),
    .A2(_13879_),
    .B1(_13885_),
    .Y(_13890_));
 sky130_fd_sc_hd__nand2_2 _23813_ (.A(_13886_),
    .B(_13889_),
    .Y(_13891_));
 sky130_fd_sc_hd__nor4_1 _23814_ (.A(_12124_),
    .B(_12127_),
    .C(_12561_),
    .D(_12563_),
    .Y(_13892_));
 sky130_fd_sc_hd__nand3_1 _23815_ (.A(_12562_),
    .B(_12564_),
    .C(_12129_),
    .Y(_13893_));
 sky130_fd_sc_hd__a211oi_2 _23816_ (.A1(_13004_),
    .A2(_13021_),
    .B1(_13893_),
    .C1(_13024_),
    .Y(_13894_));
 sky130_fd_sc_hd__nand3_1 _23817_ (.A(_13455_),
    .B(_13892_),
    .C(_13026_),
    .Y(_13895_));
 sky130_fd_sc_hd__a32oi_1 _23818_ (.A1(_07936_),
    .A2(_13450_),
    .A3(_13451_),
    .B1(_13894_),
    .B2(_13455_),
    .Y(_13896_));
 sky130_fd_sc_hd__o211a_1 _23819_ (.A1(_13460_),
    .A2(_13454_),
    .B1(_13456_),
    .C1(_13895_),
    .X(_13897_));
 sky130_fd_sc_hd__o211ai_4 _23820_ (.A1(_13460_),
    .A2(_13454_),
    .B1(_13456_),
    .C1(_13895_),
    .Y(_13899_));
 sky130_fd_sc_hd__o2111a_1 _23821_ (.A1(_12135_),
    .A2(_12138_),
    .B1(_13023_),
    .C1(_13892_),
    .D1(_13025_),
    .X(_13900_));
 sky130_fd_sc_hd__o211ai_2 _23822_ (.A1(_12135_),
    .A2(_12138_),
    .B1(_13894_),
    .C1(_13456_),
    .Y(_13901_));
 sky130_fd_sc_hd__nand3_4 _23823_ (.A(_13900_),
    .B(_13456_),
    .C(_13455_),
    .Y(_13902_));
 sky130_fd_sc_hd__a2bb2oi_1 _23824_ (.A1_N(_13454_),
    .A2_N(_13901_),
    .B1(_13462_),
    .B2(_13896_),
    .Y(_13903_));
 sky130_fd_sc_hd__o21ai_2 _23825_ (.A1(_13454_),
    .A2(_13901_),
    .B1(_13899_),
    .Y(_13904_));
 sky130_fd_sc_hd__a21oi_2 _23826_ (.A1(_13899_),
    .A2(_13902_),
    .B1(_13891_),
    .Y(_13905_));
 sky130_fd_sc_hd__a31o_1 _23827_ (.A1(_13891_),
    .A2(_13899_),
    .A3(_13902_),
    .B1(_04040_),
    .X(_13906_));
 sky130_fd_sc_hd__nand3_1 _23828_ (.A(_13886_),
    .B(_13889_),
    .C(_13902_),
    .Y(_13907_));
 sky130_fd_sc_hd__nand3_2 _23829_ (.A(_13890_),
    .B(_13899_),
    .C(_13902_),
    .Y(_13908_));
 sky130_fd_sc_hd__a22o_1 _23830_ (.A1(_13886_),
    .A2(_13889_),
    .B1(_13899_),
    .B2(_13902_),
    .X(_13910_));
 sky130_fd_sc_hd__o211a_1 _23831_ (.A1(net278),
    .A2(_13868_),
    .B1(_13878_),
    .C1(_04040_),
    .X(_13911_));
 sky130_fd_sc_hd__a311o_1 _23832_ (.A1(_13877_),
    .A2(net278),
    .A3(_13875_),
    .B1(net277),
    .C1(_13869_),
    .X(_13912_));
 sky130_fd_sc_hd__o221ai_4 _23833_ (.A1(net302),
    .A2(_04019_),
    .B1(_13890_),
    .B2(_13903_),
    .C1(_13908_),
    .Y(_13913_));
 sky130_fd_sc_hd__o221a_2 _23834_ (.A1(net277),
    .A2(_13883_),
    .B1(_13905_),
    .B2(_13906_),
    .C1(_05234_),
    .X(_13914_));
 sky130_fd_sc_hd__a211o_2 _23835_ (.A1(_13912_),
    .A2(_13913_),
    .B1(net296),
    .C1(_05232_),
    .X(_13915_));
 sky130_fd_sc_hd__a311oi_4 _23836_ (.A1(_13910_),
    .A2(net277),
    .A3(_13908_),
    .B1(_13911_),
    .C1(_07936_),
    .Y(_13916_));
 sky130_fd_sc_hd__nand3_4 _23837_ (.A(_13913_),
    .B(_07935_),
    .C(_13912_),
    .Y(_13917_));
 sky130_fd_sc_hd__o221ai_4 _23838_ (.A1(net277),
    .A2(_13883_),
    .B1(_13905_),
    .B2(_13906_),
    .C1(_07936_),
    .Y(_13918_));
 sky130_fd_sc_hd__a21oi_1 _23839_ (.A1(_13039_),
    .A2(_13466_),
    .B1(_13472_),
    .Y(_13919_));
 sky130_fd_sc_hd__a31o_1 _23840_ (.A1(_13039_),
    .A2(_13466_),
    .A3(_13471_),
    .B1(_13472_),
    .X(_13921_));
 sky130_fd_sc_hd__a31oi_4 _23841_ (.A1(_13039_),
    .A2(_13466_),
    .A3(_13471_),
    .B1(_13472_),
    .Y(_13922_));
 sky130_fd_sc_hd__o2bb2ai_4 _23842_ (.A1_N(_13917_),
    .A2_N(_13918_),
    .B1(_13919_),
    .B2(_13469_),
    .Y(_13923_));
 sky130_fd_sc_hd__nand3_4 _23843_ (.A(_13921_),
    .B(_13918_),
    .C(_13917_),
    .Y(_13924_));
 sky130_fd_sc_hd__and3_1 _23844_ (.A(_13923_),
    .B(_13924_),
    .C(net272),
    .X(_13925_));
 sky130_fd_sc_hd__nand3_2 _23845_ (.A(_13923_),
    .B(_13924_),
    .C(net272),
    .Y(_13926_));
 sky130_fd_sc_hd__a31oi_4 _23846_ (.A1(_13923_),
    .A2(_13924_),
    .A3(net272),
    .B1(_13914_),
    .Y(_13927_));
 sky130_fd_sc_hd__inv_2 _23847_ (.A(_13927_),
    .Y(_13928_));
 sky130_fd_sc_hd__o221ai_4 _23848_ (.A1(net227),
    .A2(_13052_),
    .B1(_13490_),
    .B2(_13068_),
    .C1(_13486_),
    .Y(_13929_));
 sky130_fd_sc_hd__o21ai_1 _23849_ (.A1(net222),
    .A2(_13483_),
    .B1(_13491_),
    .Y(_13930_));
 sky130_fd_sc_hd__a311oi_4 _23850_ (.A1(_13923_),
    .A2(_13924_),
    .A3(net272),
    .B1(net202),
    .C1(_13914_),
    .Y(_13932_));
 sky130_fd_sc_hd__nand3_2 _23851_ (.A(_13926_),
    .B(_07564_),
    .C(_13915_),
    .Y(_13933_));
 sky130_fd_sc_hd__a22oi_4 _23852_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_13915_),
    .B2(_13926_),
    .Y(_13934_));
 sky130_fd_sc_hd__a22o_1 _23853_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_13915_),
    .B2(_13926_),
    .X(_13935_));
 sky130_fd_sc_hd__nor2_1 _23854_ (.A(_13932_),
    .B(_13934_),
    .Y(_13936_));
 sky130_fd_sc_hd__o2111ai_1 _23855_ (.A1(_13484_),
    .A2(net224),
    .B1(_13933_),
    .C1(_13930_),
    .D1(_13935_),
    .Y(_13937_));
 sky130_fd_sc_hd__o221ai_2 _23856_ (.A1(net222),
    .A2(_13483_),
    .B1(_13932_),
    .B2(_13934_),
    .C1(_13929_),
    .Y(_13938_));
 sky130_fd_sc_hd__o211ai_2 _23857_ (.A1(net270),
    .A2(net268),
    .B1(_13937_),
    .C1(_13938_),
    .Y(_13939_));
 sky130_fd_sc_hd__o221ai_4 _23858_ (.A1(_13483_),
    .A2(net222),
    .B1(_07564_),
    .B2(_13927_),
    .C1(_13929_),
    .Y(_13940_));
 sky130_fd_sc_hd__o2bb2ai_1 _23859_ (.A1_N(_13488_),
    .A2_N(_13929_),
    .B1(_13932_),
    .B2(_13934_),
    .Y(_13941_));
 sky130_fd_sc_hd__o221ai_4 _23860_ (.A1(net270),
    .A2(net268),
    .B1(_13932_),
    .B2(_13940_),
    .C1(_13941_),
    .Y(_13943_));
 sky130_fd_sc_hd__o31a_1 _23861_ (.A1(net245),
    .A2(_13914_),
    .A3(_13925_),
    .B1(_13939_),
    .X(_13944_));
 sky130_fd_sc_hd__o31a_2 _23862_ (.A1(net270),
    .A2(net268),
    .A3(_13927_),
    .B1(_13943_),
    .X(_13945_));
 sky130_fd_sc_hd__o311a_2 _23863_ (.A1(net270),
    .A2(net268),
    .A3(_13927_),
    .B1(_13943_),
    .C1(_05754_),
    .X(_13946_));
 sky130_fd_sc_hd__o211ai_4 _23864_ (.A1(_13928_),
    .A2(net245),
    .B1(net222),
    .C1(_13939_),
    .Y(_13947_));
 sky130_fd_sc_hd__o211ai_4 _23865_ (.A1(net245),
    .A2(_13927_),
    .B1(_07246_),
    .C1(_13943_),
    .Y(_13948_));
 sky130_fd_sc_hd__nand2_1 _23866_ (.A(_13947_),
    .B(_13948_),
    .Y(_13949_));
 sky130_fd_sc_hd__a22o_1 _23867_ (.A1(net225),
    .A2(_13502_),
    .B1(_13517_),
    .B2(_13519_),
    .X(_13950_));
 sky130_fd_sc_hd__o211ai_4 _23868_ (.A1(_13507_),
    .A2(_13499_),
    .B1(_13519_),
    .C1(_13517_),
    .Y(_13951_));
 sky130_fd_sc_hd__o2111ai_4 _23869_ (.A1(net227),
    .A2(_13501_),
    .B1(_13947_),
    .C1(_13948_),
    .D1(_13951_),
    .Y(_13952_));
 sky130_fd_sc_hd__o221ai_4 _23870_ (.A1(_13507_),
    .A2(_13499_),
    .B1(_13504_),
    .B2(_13520_),
    .C1(_13949_),
    .Y(_13954_));
 sky130_fd_sc_hd__o211ai_2 _23871_ (.A1(_05750_),
    .A2(net264),
    .B1(_13952_),
    .C1(_13954_),
    .Y(_13955_));
 sky130_fd_sc_hd__or3_2 _23872_ (.A(_05750_),
    .B(net264),
    .C(_13945_),
    .X(_13956_));
 sky130_fd_sc_hd__o221ai_2 _23873_ (.A1(net227),
    .A2(_13501_),
    .B1(_13511_),
    .B2(_13521_),
    .C1(_13949_),
    .Y(_13957_));
 sky130_fd_sc_hd__o2111ai_1 _23874_ (.A1(net225),
    .A2(_13502_),
    .B1(_13947_),
    .C1(_13948_),
    .D1(_13950_),
    .Y(_13958_));
 sky130_fd_sc_hd__nand3_1 _23875_ (.A(_13958_),
    .B(net243),
    .C(_13957_),
    .Y(_13959_));
 sky130_fd_sc_hd__a31o_4 _23876_ (.A1(_13954_),
    .A2(net243),
    .A3(_13952_),
    .B1(_13946_),
    .X(_13960_));
 sky130_fd_sc_hd__inv_2 _23877_ (.A(_13960_),
    .Y(_13961_));
 sky130_fd_sc_hd__a311o_1 _23878_ (.A1(_13954_),
    .A2(net243),
    .A3(_13952_),
    .B1(net240),
    .C1(_13946_),
    .X(_13962_));
 sky130_fd_sc_hd__nand4_1 _23879_ (.A(_12201_),
    .B(_12203_),
    .C(_12635_),
    .D(_12638_),
    .Y(_13963_));
 sky130_fd_sc_hd__nor3_1 _23880_ (.A(_13107_),
    .B(_13963_),
    .C(_13110_),
    .Y(_13965_));
 sky130_fd_sc_hd__nand2_1 _23881_ (.A(_13535_),
    .B(_13965_),
    .Y(_13966_));
 sky130_fd_sc_hd__o211a_2 _23882_ (.A1(_13541_),
    .A2(_13534_),
    .B1(_13537_),
    .C1(_13966_),
    .X(_13967_));
 sky130_fd_sc_hd__o211ai_4 _23883_ (.A1(_13541_),
    .A2(_13534_),
    .B1(_13537_),
    .C1(_13966_),
    .Y(_13968_));
 sky130_fd_sc_hd__nand4_4 _23884_ (.A(_13535_),
    .B(_13537_),
    .C(_13965_),
    .D(_12216_),
    .Y(_13969_));
 sky130_fd_sc_hd__inv_2 _23885_ (.A(_13969_),
    .Y(_13970_));
 sky130_fd_sc_hd__a31o_1 _23886_ (.A1(_13537_),
    .A2(_13545_),
    .A3(_13966_),
    .B1(_13970_),
    .X(_13971_));
 sky130_fd_sc_hd__a311oi_4 _23887_ (.A1(_13954_),
    .A2(net243),
    .A3(_13952_),
    .B1(net227),
    .C1(_13946_),
    .Y(_13972_));
 sky130_fd_sc_hd__o211ai_4 _23888_ (.A1(net243),
    .A2(_13944_),
    .B1(_13955_),
    .C1(net225),
    .Y(_13973_));
 sky130_fd_sc_hd__a31oi_1 _23889_ (.A1(_13958_),
    .A2(net243),
    .A3(_13957_),
    .B1(net225),
    .Y(_13974_));
 sky130_fd_sc_hd__and3_1 _23890_ (.A(_13959_),
    .B(net227),
    .C(_13956_),
    .X(_13976_));
 sky130_fd_sc_hd__nand3_4 _23891_ (.A(_13959_),
    .B(net227),
    .C(_13956_),
    .Y(_13977_));
 sky130_fd_sc_hd__a21oi_1 _23892_ (.A1(_13974_),
    .A2(_13956_),
    .B1(_13972_),
    .Y(_13978_));
 sky130_fd_sc_hd__a21oi_2 _23893_ (.A1(_13968_),
    .A2(_13969_),
    .B1(_13978_),
    .Y(_13979_));
 sky130_fd_sc_hd__o2bb2ai_4 _23894_ (.A1_N(_13968_),
    .A2_N(_13969_),
    .B1(_13972_),
    .B2(_13976_),
    .Y(_13980_));
 sky130_fd_sc_hd__nand3_1 _23895_ (.A(_13969_),
    .B(_13973_),
    .C(_13977_),
    .Y(_13981_));
 sky130_fd_sc_hd__a41oi_4 _23896_ (.A1(_13968_),
    .A2(_13969_),
    .A3(_13973_),
    .A4(_13977_),
    .B1(_05995_),
    .Y(_13982_));
 sky130_fd_sc_hd__o22ai_4 _23897_ (.A1(net260),
    .A2(net258),
    .B1(_13981_),
    .B2(_13967_),
    .Y(_13983_));
 sky130_fd_sc_hd__nand2_1 _23898_ (.A(_13982_),
    .B(_13980_),
    .Y(_13984_));
 sky130_fd_sc_hd__a22oi_4 _23899_ (.A1(_05995_),
    .A2(_13961_),
    .B1(_13982_),
    .B2(_13980_),
    .Y(_13985_));
 sky130_fd_sc_hd__o22ai_2 _23900_ (.A1(net240),
    .A2(_13960_),
    .B1(_13979_),
    .B2(_13983_),
    .Y(_13987_));
 sky130_fd_sc_hd__a21oi_2 _23901_ (.A1(_13962_),
    .A2(_13984_),
    .B1(net214),
    .Y(_13988_));
 sky130_fd_sc_hd__or3_1 _23902_ (.A(net239),
    .B(_06292_),
    .C(_13985_),
    .X(_13989_));
 sky130_fd_sc_hd__a221oi_4 _23903_ (.A1(_05995_),
    .A2(_13961_),
    .B1(_13982_),
    .B2(_13980_),
    .C1(net233),
    .Y(_13990_));
 sky130_fd_sc_hd__o221ai_4 _23904_ (.A1(net240),
    .A2(_13960_),
    .B1(_13979_),
    .B2(_13983_),
    .C1(net234),
    .Y(_13991_));
 sky130_fd_sc_hd__a2bb2oi_1 _23905_ (.A1_N(_06622_),
    .A2_N(_06624_),
    .B1(_13962_),
    .B2(_13984_),
    .Y(_13992_));
 sky130_fd_sc_hd__o21ai_4 _23906_ (.A1(_06622_),
    .A2(_06624_),
    .B1(_13987_),
    .Y(_13993_));
 sky130_fd_sc_hd__a21o_1 _23907_ (.A1(_13552_),
    .A2(_13554_),
    .B1(_13555_),
    .X(_13994_));
 sky130_fd_sc_hd__a21oi_2 _23908_ (.A1(_13552_),
    .A2(_13554_),
    .B1(_13555_),
    .Y(_13995_));
 sky130_fd_sc_hd__a21oi_2 _23909_ (.A1(_13991_),
    .A2(_13993_),
    .B1(_13994_),
    .Y(_13996_));
 sky130_fd_sc_hd__o21ai_4 _23910_ (.A1(_13990_),
    .A2(_13992_),
    .B1(_13995_),
    .Y(_13998_));
 sky130_fd_sc_hd__o21ai_1 _23911_ (.A1(net235),
    .A2(_13985_),
    .B1(_13994_),
    .Y(_13999_));
 sky130_fd_sc_hd__nand3_2 _23912_ (.A(_13991_),
    .B(_13993_),
    .C(_13994_),
    .Y(_14000_));
 sky130_fd_sc_hd__o22ai_4 _23913_ (.A1(net239),
    .A2(_06292_),
    .B1(_13990_),
    .B2(_13999_),
    .Y(_14001_));
 sky130_fd_sc_hd__nand3_1 _23914_ (.A(_13998_),
    .B(_14000_),
    .C(net213),
    .Y(_14002_));
 sky130_fd_sc_hd__a31oi_4 _23915_ (.A1(_13998_),
    .A2(_14000_),
    .A3(net214),
    .B1(_13988_),
    .Y(_14003_));
 sky130_fd_sc_hd__o22ai_4 _23916_ (.A1(net213),
    .A2(_13985_),
    .B1(_13996_),
    .B2(_14001_),
    .Y(_14004_));
 sky130_fd_sc_hd__o311a_1 _23917_ (.A1(_05765_),
    .A2(_13142_),
    .A3(_05766_),
    .B1(_13571_),
    .C1(_13158_),
    .X(_14005_));
 sky130_fd_sc_hd__a21oi_1 _23918_ (.A1(_13143_),
    .A2(_13158_),
    .B1(_13567_),
    .Y(_14006_));
 sky130_fd_sc_hd__a31oi_2 _23919_ (.A1(_13143_),
    .A2(_13158_),
    .A3(_13571_),
    .B1(_13567_),
    .Y(_14007_));
 sky130_fd_sc_hd__a311oi_4 _23920_ (.A1(_13998_),
    .A2(_14000_),
    .A3(net214),
    .B1(net252),
    .C1(_13988_),
    .Y(_14009_));
 sky130_fd_sc_hd__o221ai_4 _23921_ (.A1(net213),
    .A2(_13985_),
    .B1(_13996_),
    .B2(_14001_),
    .C1(_06314_),
    .Y(_14010_));
 sky130_fd_sc_hd__a2bb2oi_2 _23922_ (.A1_N(net284),
    .A2_N(net282),
    .B1(_13989_),
    .B2(_14002_),
    .Y(_14011_));
 sky130_fd_sc_hd__o21ai_1 _23923_ (.A1(net284),
    .A2(net282),
    .B1(_14004_),
    .Y(_14012_));
 sky130_fd_sc_hd__nor2_1 _23924_ (.A(_14009_),
    .B(_14011_),
    .Y(_14013_));
 sky130_fd_sc_hd__o211ai_1 _23925_ (.A1(_13567_),
    .A2(_14005_),
    .B1(_14010_),
    .C1(_14012_),
    .Y(_14014_));
 sky130_fd_sc_hd__o22ai_1 _23926_ (.A1(_13570_),
    .A2(_14006_),
    .B1(_14009_),
    .B2(_14011_),
    .Y(_14015_));
 sky130_fd_sc_hd__nand3_1 _23927_ (.A(_14014_),
    .B(_14015_),
    .C(net210),
    .Y(_14016_));
 sky130_fd_sc_hd__or3_1 _23928_ (.A(net238),
    .B(_06610_),
    .C(_14003_),
    .X(_14017_));
 sky130_fd_sc_hd__o21ai_1 _23929_ (.A1(_06314_),
    .A2(_14003_),
    .B1(_14007_),
    .Y(_14018_));
 sky130_fd_sc_hd__o22ai_2 _23930_ (.A1(_13567_),
    .A2(_14005_),
    .B1(_14009_),
    .B2(_14011_),
    .Y(_14020_));
 sky130_fd_sc_hd__o221ai_4 _23931_ (.A1(net238),
    .A2(_06610_),
    .B1(_14009_),
    .B2(_14018_),
    .C1(_14020_),
    .Y(_14021_));
 sky130_fd_sc_hd__o21ai_4 _23932_ (.A1(net210),
    .A2(_14003_),
    .B1(_14021_),
    .Y(_14022_));
 sky130_fd_sc_hd__o211a_1 _23933_ (.A1(_14004_),
    .A2(net210),
    .B1(_06014_),
    .C1(_14016_),
    .X(_14023_));
 sky130_fd_sc_hd__o211ai_4 _23934_ (.A1(_14004_),
    .A2(net210),
    .B1(_06014_),
    .C1(_14016_),
    .Y(_14024_));
 sky130_fd_sc_hd__o221a_2 _23935_ (.A1(_06011_),
    .A2(_06012_),
    .B1(net210),
    .B2(_14003_),
    .C1(_14021_),
    .X(_14025_));
 sky130_fd_sc_hd__o221ai_4 _23936_ (.A1(_06011_),
    .A2(_06012_),
    .B1(net210),
    .B2(_14003_),
    .C1(_14021_),
    .Y(_14026_));
 sky130_fd_sc_hd__nand2_1 _23937_ (.A(_14024_),
    .B(_14026_),
    .Y(_14027_));
 sky130_fd_sc_hd__o22ai_2 _23938_ (.A1(net263),
    .A2(_13583_),
    .B1(_13608_),
    .B2(_13596_),
    .Y(_14028_));
 sky130_fd_sc_hd__and4_1 _23939_ (.A(_13586_),
    .B(_13609_),
    .C(_14024_),
    .D(_14026_),
    .X(_14029_));
 sky130_fd_sc_hd__o2bb2ai_2 _23940_ (.A1_N(_14028_),
    .A2_N(_14027_),
    .B1(net228),
    .B2(net231),
    .Y(_14031_));
 sky130_fd_sc_hd__and3_1 _23941_ (.A(_14022_),
    .B(_06902_),
    .C(_06900_),
    .X(_14032_));
 sky130_fd_sc_hd__a211o_1 _23942_ (.A1(_14017_),
    .A2(_14021_),
    .B1(net231),
    .C1(net228),
    .X(_14033_));
 sky130_fd_sc_hd__o221ai_2 _23943_ (.A1(net263),
    .A2(_13583_),
    .B1(_13596_),
    .B2(_13608_),
    .C1(_14027_),
    .Y(_14034_));
 sky130_fd_sc_hd__nand3_1 _23944_ (.A(_14028_),
    .B(_14026_),
    .C(_14024_),
    .Y(_14035_));
 sky130_fd_sc_hd__nand3_1 _23945_ (.A(_14034_),
    .B(_14035_),
    .C(net208),
    .Y(_14036_));
 sky130_fd_sc_hd__a31o_2 _23946_ (.A1(_14034_),
    .A2(_14035_),
    .A3(net208),
    .B1(_14032_),
    .X(_14037_));
 sky130_fd_sc_hd__o221a_2 _23947_ (.A1(net208),
    .A2(_14022_),
    .B1(_14029_),
    .B2(_14031_),
    .C1(_05768_),
    .X(_14038_));
 sky130_fd_sc_hd__o221ai_4 _23948_ (.A1(net208),
    .A2(_14022_),
    .B1(_14029_),
    .B2(_14031_),
    .C1(_05768_),
    .Y(_14039_));
 sky130_fd_sc_hd__nand3_4 _23949_ (.A(_14036_),
    .B(net263),
    .C(_14033_),
    .Y(_14040_));
 sky130_fd_sc_hd__nand2_1 _23950_ (.A(_14039_),
    .B(_14040_),
    .Y(_14042_));
 sky130_fd_sc_hd__nand4_1 _23951_ (.A(_12274_),
    .B(_12277_),
    .C(_12707_),
    .D(_12709_),
    .Y(_14043_));
 sky130_fd_sc_hd__a211oi_2 _23952_ (.A1(_13162_),
    .A2(_13184_),
    .B1(_14043_),
    .C1(_13188_),
    .Y(_14044_));
 sky130_fd_sc_hd__nand2_1 _23953_ (.A(_13617_),
    .B(_14044_),
    .Y(_14045_));
 sky130_fd_sc_hd__o211ai_4 _23954_ (.A1(_13622_),
    .A2(_13616_),
    .B1(_13618_),
    .C1(_14045_),
    .Y(_14046_));
 sky130_fd_sc_hd__nand4_4 _23955_ (.A(_14044_),
    .B(_13618_),
    .C(_13617_),
    .D(_11959_),
    .Y(_14047_));
 sky130_fd_sc_hd__nand2_1 _23956_ (.A(_14046_),
    .B(_14047_),
    .Y(_14048_));
 sky130_fd_sc_hd__a21oi_2 _23957_ (.A1(_14046_),
    .A2(_14047_),
    .B1(_14042_),
    .Y(_14049_));
 sky130_fd_sc_hd__a31o_1 _23958_ (.A1(_14042_),
    .A2(_14046_),
    .A3(_14047_),
    .B1(_07232_),
    .X(_14050_));
 sky130_fd_sc_hd__a211o_2 _23959_ (.A1(_14033_),
    .A2(_14036_),
    .B1(net207),
    .C1(net206),
    .X(_14051_));
 sky130_fd_sc_hd__a22oi_1 _23960_ (.A1(_14039_),
    .A2(_14040_),
    .B1(_14046_),
    .B2(_14047_),
    .Y(_14053_));
 sky130_fd_sc_hd__a22o_1 _23961_ (.A1(_14039_),
    .A2(_14040_),
    .B1(_14046_),
    .B2(_14047_),
    .X(_14054_));
 sky130_fd_sc_hd__o211ai_4 _23962_ (.A1(_14037_),
    .A2(_05768_),
    .B1(_14047_),
    .C1(_14046_),
    .Y(_14055_));
 sky130_fd_sc_hd__o2111a_1 _23963_ (.A1(_05768_),
    .A2(_14037_),
    .B1(_14039_),
    .C1(_14046_),
    .D1(_14047_),
    .X(_14056_));
 sky130_fd_sc_hd__o221ai_4 _23964_ (.A1(_07227_),
    .A2(net206),
    .B1(_14038_),
    .B2(_14055_),
    .C1(_14054_),
    .Y(_14057_));
 sky130_fd_sc_hd__o31a_1 _23965_ (.A1(_07232_),
    .A2(_14053_),
    .A3(_14056_),
    .B1(_14051_),
    .X(_14058_));
 sky130_fd_sc_hd__o221a_2 _23966_ (.A1(net185),
    .A2(_14037_),
    .B1(_14049_),
    .B2(_14050_),
    .C1(_07550_),
    .X(_14059_));
 sky130_fd_sc_hd__a211o_1 _23967_ (.A1(_14051_),
    .A2(_14057_),
    .B1(_07544_),
    .C1(_07546_),
    .X(_14060_));
 sky130_fd_sc_hd__o311a_1 _23968_ (.A1(_07232_),
    .A2(_14053_),
    .A3(_14056_),
    .B1(_14051_),
    .C1(_05507_),
    .X(_14061_));
 sky130_fd_sc_hd__nand3_4 _23969_ (.A(_14057_),
    .B(_05507_),
    .C(_14051_),
    .Y(_14062_));
 sky130_fd_sc_hd__o221ai_4 _23970_ (.A1(net185),
    .A2(_14037_),
    .B1(_14049_),
    .B2(_14050_),
    .C1(net292),
    .Y(_14064_));
 sky130_fd_sc_hd__o211a_1 _23971_ (.A1(_13206_),
    .A2(_13202_),
    .B1(_13201_),
    .C1(_13641_),
    .X(_14065_));
 sky130_fd_sc_hd__o311a_1 _23972_ (.A1(_12720_),
    .A2(_12733_),
    .A3(_13200_),
    .B1(_13203_),
    .C1(_13639_),
    .X(_14066_));
 sky130_fd_sc_hd__a21oi_2 _23973_ (.A1(_13639_),
    .A2(_13636_),
    .B1(_13640_),
    .Y(_14067_));
 sky130_fd_sc_hd__a21boi_1 _23974_ (.A1(_14062_),
    .A2(_14064_),
    .B1_N(_14067_),
    .Y(_14068_));
 sky130_fd_sc_hd__o2bb2ai_4 _23975_ (.A1_N(_14062_),
    .A2_N(_14064_),
    .B1(_14065_),
    .B2(_13638_),
    .Y(_14069_));
 sky130_fd_sc_hd__o211a_1 _23976_ (.A1(_13640_),
    .A2(_14066_),
    .B1(_14064_),
    .C1(_14062_),
    .X(_14070_));
 sky130_fd_sc_hd__o211ai_4 _23977_ (.A1(_13640_),
    .A2(_14066_),
    .B1(_14064_),
    .C1(_14062_),
    .Y(_14071_));
 sky130_fd_sc_hd__nand3_2 _23978_ (.A(_14069_),
    .B(_14071_),
    .C(net163),
    .Y(_14072_));
 sky130_fd_sc_hd__nand2_1 _23979_ (.A(_07550_),
    .B(_14058_),
    .Y(_14073_));
 sky130_fd_sc_hd__o22ai_1 _23980_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_14068_),
    .B2(_14070_),
    .Y(_14075_));
 sky130_fd_sc_hd__a31oi_2 _23981_ (.A1(_14069_),
    .A2(_14071_),
    .A3(net163),
    .B1(_14059_),
    .Y(_14076_));
 sky130_fd_sc_hd__a31o_1 _23982_ (.A1(_14069_),
    .A2(_14071_),
    .A3(net163),
    .B1(_14059_),
    .X(_14077_));
 sky130_fd_sc_hd__o311a_2 _23983_ (.A1(_12742_),
    .A2(_13220_),
    .A3(_13222_),
    .B1(_13652_),
    .C1(_13219_),
    .X(_14078_));
 sky130_fd_sc_hd__a221oi_2 _23984_ (.A1(_02137_),
    .A2(_13215_),
    .B1(_13650_),
    .B2(_04227_),
    .C1(_13655_),
    .Y(_14079_));
 sky130_fd_sc_hd__nand2_1 _23985_ (.A(_13654_),
    .B(_13656_),
    .Y(_14080_));
 sky130_fd_sc_hd__o21ai_1 _23986_ (.A1(_04227_),
    .A2(_13650_),
    .B1(_14080_),
    .Y(_14081_));
 sky130_fd_sc_hd__a311oi_4 _23987_ (.A1(_14069_),
    .A2(_14071_),
    .A3(net163),
    .B1(_14059_),
    .C1(net294),
    .Y(_14082_));
 sky130_fd_sc_hd__o211ai_2 _23988_ (.A1(net163),
    .A2(_14058_),
    .B1(net295),
    .C1(_14072_),
    .Y(_14083_));
 sky130_fd_sc_hd__a2bb2oi_4 _23989_ (.A1_N(net318),
    .A2_N(net316),
    .B1(_14060_),
    .B2(_14072_),
    .Y(_14084_));
 sky130_fd_sc_hd__o211ai_2 _23990_ (.A1(net318),
    .A2(net316),
    .B1(_14073_),
    .C1(_14075_),
    .Y(_14086_));
 sky130_fd_sc_hd__o211ai_1 _23991_ (.A1(_13653_),
    .A2(_14078_),
    .B1(_14083_),
    .C1(_14086_),
    .Y(_14087_));
 sky130_fd_sc_hd__o22ai_1 _23992_ (.A1(_13651_),
    .A2(_14079_),
    .B1(_14082_),
    .B2(_14084_),
    .Y(_14088_));
 sky130_fd_sc_hd__o211ai_2 _23993_ (.A1(net183),
    .A2(net182),
    .B1(_14087_),
    .C1(_14088_),
    .Y(_14089_));
 sky130_fd_sc_hd__and3_1 _23994_ (.A(_07917_),
    .B(_14073_),
    .C(_14075_),
    .X(_14090_));
 sky130_fd_sc_hd__nand3_2 _23995_ (.A(_14086_),
    .B(_14081_),
    .C(_14083_),
    .Y(_14091_));
 sky130_fd_sc_hd__o22ai_4 _23996_ (.A1(_13653_),
    .A2(_14078_),
    .B1(_14082_),
    .B2(_14084_),
    .Y(_14092_));
 sky130_fd_sc_hd__o211ai_2 _23997_ (.A1(net183),
    .A2(net182),
    .B1(_14091_),
    .C1(_14092_),
    .Y(_14093_));
 sky130_fd_sc_hd__a31oi_4 _23998_ (.A1(_14092_),
    .A2(net161),
    .A3(_14091_),
    .B1(_14090_),
    .Y(_14094_));
 sky130_fd_sc_hd__o211a_1 _23999_ (.A1(_14077_),
    .A2(net161),
    .B1(_04238_),
    .C1(_14089_),
    .X(_14095_));
 sky130_fd_sc_hd__o211ai_4 _24000_ (.A1(_14077_),
    .A2(net161),
    .B1(_04238_),
    .C1(_14089_),
    .Y(_14097_));
 sky130_fd_sc_hd__o211a_2 _24001_ (.A1(net161),
    .A2(_14076_),
    .B1(_04227_),
    .C1(_14093_),
    .X(_14098_));
 sky130_fd_sc_hd__o211ai_2 _24002_ (.A1(net161),
    .A2(_14076_),
    .B1(_04227_),
    .C1(_14093_),
    .Y(_14099_));
 sky130_fd_sc_hd__a21oi_1 _24003_ (.A1(_13675_),
    .A2(_13677_),
    .B1(_13664_),
    .Y(_14100_));
 sky130_fd_sc_hd__a31o_1 _24004_ (.A1(_13667_),
    .A2(_13675_),
    .A3(_13677_),
    .B1(_13664_),
    .X(_14101_));
 sky130_fd_sc_hd__a31oi_2 _24005_ (.A1(_13667_),
    .A2(_13675_),
    .A3(_13677_),
    .B1(_13664_),
    .Y(_14102_));
 sky130_fd_sc_hd__o2bb2ai_1 _24006_ (.A1_N(_14097_),
    .A2_N(_14099_),
    .B1(_14100_),
    .B2(_13666_),
    .Y(_14103_));
 sky130_fd_sc_hd__nand3_1 _24007_ (.A(_14101_),
    .B(_14099_),
    .C(_14097_),
    .Y(_14104_));
 sky130_fd_sc_hd__nand3_4 _24008_ (.A(_14103_),
    .B(_14104_),
    .C(_08300_),
    .Y(_14105_));
 sky130_fd_sc_hd__or3_2 _24009_ (.A(net180),
    .B(_08298_),
    .C(_14094_),
    .X(_14106_));
 sky130_fd_sc_hd__o31a_1 _24010_ (.A1(net180),
    .A2(_08298_),
    .A3(_14094_),
    .B1(_14105_),
    .X(_14108_));
 sky130_fd_sc_hd__inv_2 _24011_ (.A(_14108_),
    .Y(_14109_));
 sky130_fd_sc_hd__a22oi_2 _24012_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_14105_),
    .B2(_14106_),
    .Y(_14110_));
 sky130_fd_sc_hd__a22o_1 _24013_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_14105_),
    .B2(_14106_),
    .X(_14111_));
 sky130_fd_sc_hd__o211a_2 _24014_ (.A1(_08300_),
    .A2(_14094_),
    .B1(_02137_),
    .C1(_14105_),
    .X(_14112_));
 sky130_fd_sc_hd__o211ai_2 _24015_ (.A1(_08300_),
    .A2(_14094_),
    .B1(_02137_),
    .C1(_14105_),
    .Y(_14113_));
 sky130_fd_sc_hd__o22a_1 _24016_ (.A1(_13692_),
    .A2(_13686_),
    .B1(_13697_),
    .B2(_13694_),
    .X(_14114_));
 sky130_fd_sc_hd__o22ai_4 _24017_ (.A1(_13692_),
    .A2(_13686_),
    .B1(_13697_),
    .B2(_13694_),
    .Y(_14115_));
 sky130_fd_sc_hd__nand3_1 _24018_ (.A(_14111_),
    .B(_14113_),
    .C(_14115_),
    .Y(_14116_));
 sky130_fd_sc_hd__o21ai_1 _24019_ (.A1(_14110_),
    .A2(_14112_),
    .B1(_14114_),
    .Y(_14117_));
 sky130_fd_sc_hd__nand3_2 _24020_ (.A(_14117_),
    .B(_08714_),
    .C(_14116_),
    .Y(_14119_));
 sky130_fd_sc_hd__a21oi_1 _24021_ (.A1(_14105_),
    .A2(_14106_),
    .B1(_08714_),
    .Y(_14120_));
 sky130_fd_sc_hd__a22o_1 _24022_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_14105_),
    .B2(_14106_),
    .X(_14121_));
 sky130_fd_sc_hd__o21ai_2 _24023_ (.A1(_14110_),
    .A2(_14112_),
    .B1(_14115_),
    .Y(_14122_));
 sky130_fd_sc_hd__nand3_1 _24024_ (.A(_14111_),
    .B(_14114_),
    .C(_14113_),
    .Y(_14123_));
 sky130_fd_sc_hd__nand3_1 _24025_ (.A(_14122_),
    .B(_14123_),
    .C(_08714_),
    .Y(_14124_));
 sky130_fd_sc_hd__a31o_1 _24026_ (.A1(_14122_),
    .A2(_14123_),
    .A3(_08714_),
    .B1(_14120_),
    .X(_14125_));
 sky130_fd_sc_hd__o311a_4 _24027_ (.A1(net158),
    .A2(_08712_),
    .A3(_14109_),
    .B1(_09124_),
    .C1(_14119_),
    .X(_14126_));
 sky130_fd_sc_hd__a211o_1 _24028_ (.A1(_14121_),
    .A2(_14124_),
    .B1(_09120_),
    .C1(_09121_),
    .X(_14127_));
 sky130_fd_sc_hd__a311oi_2 _24029_ (.A1(_14122_),
    .A2(_14123_),
    .A3(_08714_),
    .B1(_14120_),
    .C1(_00251_),
    .Y(_14128_));
 sky130_fd_sc_hd__nand3_4 _24030_ (.A(_14124_),
    .B(_00240_),
    .C(_14121_),
    .Y(_14130_));
 sky130_fd_sc_hd__o211a_2 _24031_ (.A1(_14109_),
    .A2(_08714_),
    .B1(_00251_),
    .C1(_14119_),
    .X(_14131_));
 sky130_fd_sc_hd__o211ai_4 _24032_ (.A1(_14109_),
    .A2(_08714_),
    .B1(_00251_),
    .C1(_14119_),
    .Y(_14132_));
 sky130_fd_sc_hd__o221a_1 _24033_ (.A1(_13276_),
    .A2(_13272_),
    .B1(_12888_),
    .B2(_13702_),
    .C1(_13271_),
    .X(_14133_));
 sky130_fd_sc_hd__a21oi_1 _24034_ (.A1(_12888_),
    .A2(_13702_),
    .B1(_13706_),
    .Y(_14134_));
 sky130_fd_sc_hd__a31o_1 _24035_ (.A1(_13274_),
    .A2(_13704_),
    .A3(_13708_),
    .B1(_13709_),
    .X(_14135_));
 sky130_fd_sc_hd__a21oi_2 _24036_ (.A1(_13708_),
    .A2(_13705_),
    .B1(_13709_),
    .Y(_14136_));
 sky130_fd_sc_hd__a21oi_1 _24037_ (.A1(_14130_),
    .A2(_14132_),
    .B1(_14135_),
    .Y(_14137_));
 sky130_fd_sc_hd__o2bb2ai_2 _24038_ (.A1_N(_14130_),
    .A2_N(_14132_),
    .B1(_14133_),
    .B2(_13707_),
    .Y(_14138_));
 sky130_fd_sc_hd__o211a_1 _24039_ (.A1(_13709_),
    .A2(_14134_),
    .B1(_14132_),
    .C1(_14130_),
    .X(_14139_));
 sky130_fd_sc_hd__o211ai_1 _24040_ (.A1(_13709_),
    .A2(_14134_),
    .B1(_14132_),
    .C1(_14130_),
    .Y(_14141_));
 sky130_fd_sc_hd__a31oi_2 _24041_ (.A1(_14135_),
    .A2(_14132_),
    .A3(_14130_),
    .B1(_09124_),
    .Y(_14142_));
 sky130_fd_sc_hd__nand3_1 _24042_ (.A(_09125_),
    .B(_14138_),
    .C(_14141_),
    .Y(_14143_));
 sky130_fd_sc_hd__o22ai_2 _24043_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_14137_),
    .B2(_14139_),
    .Y(_14144_));
 sky130_fd_sc_hd__o31a_2 _24044_ (.A1(_09124_),
    .A2(_14137_),
    .A3(_14139_),
    .B1(_14127_),
    .X(_14145_));
 sky130_fd_sc_hd__a311o_1 _24045_ (.A1(_09125_),
    .A2(_14138_),
    .A3(_14141_),
    .B1(net143),
    .C1(_14126_),
    .X(_14146_));
 sky130_fd_sc_hd__a21oi_2 _24046_ (.A1(_13721_),
    .A2(_11309_),
    .B1(_13729_),
    .Y(_14147_));
 sky130_fd_sc_hd__a21o_1 _24047_ (.A1(_13729_),
    .A2(_13728_),
    .B1(_13724_),
    .X(_14148_));
 sky130_fd_sc_hd__o2bb2ai_4 _24048_ (.A1_N(_14138_),
    .A2_N(_14142_),
    .B1(_12867_),
    .B2(_12877_),
    .Y(_14149_));
 sky130_fd_sc_hd__o211a_1 _24049_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_14127_),
    .C1(_14143_),
    .X(_14150_));
 sky130_fd_sc_hd__a21oi_2 _24050_ (.A1(_14127_),
    .A2(_14143_),
    .B1(_12888_),
    .Y(_14152_));
 sky130_fd_sc_hd__o211ai_4 _24051_ (.A1(_14125_),
    .A2(_09125_),
    .B1(_12899_),
    .C1(_14144_),
    .Y(_14153_));
 sky130_fd_sc_hd__o221ai_4 _24052_ (.A1(_13727_),
    .A2(_14147_),
    .B1(_14126_),
    .B2(_14149_),
    .C1(_14153_),
    .Y(_14154_));
 sky130_fd_sc_hd__o21ai_1 _24053_ (.A1(_14150_),
    .A2(_14152_),
    .B1(_14148_),
    .Y(_14155_));
 sky130_fd_sc_hd__o2111ai_4 _24054_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .C1(_14154_),
    .D1(_14155_),
    .Y(_14156_));
 sky130_fd_sc_hd__nand2_1 _24055_ (.A(_14153_),
    .B(_14148_),
    .Y(_14157_));
 sky130_fd_sc_hd__o22ai_2 _24056_ (.A1(_13727_),
    .A2(_14147_),
    .B1(_14150_),
    .B2(_14152_),
    .Y(_14158_));
 sky130_fd_sc_hd__o221ai_4 _24057_ (.A1(_09553_),
    .A2(net155),
    .B1(_14150_),
    .B2(_14157_),
    .C1(_14158_),
    .Y(_14159_));
 sky130_fd_sc_hd__o31a_2 _24058_ (.A1(_09553_),
    .A2(net155),
    .A3(_14145_),
    .B1(_14159_),
    .X(_14160_));
 sky130_fd_sc_hd__o211ai_4 _24059_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_14146_),
    .C1(_14156_),
    .Y(_14161_));
 sky130_fd_sc_hd__o211a_1 _24060_ (.A1(net143),
    .A2(_14145_),
    .B1(_11298_),
    .C1(_14159_),
    .X(_14163_));
 sky130_fd_sc_hd__o211ai_4 _24061_ (.A1(net143),
    .A2(_14145_),
    .B1(_11298_),
    .C1(_14159_),
    .Y(_14164_));
 sky130_fd_sc_hd__a2bb2oi_2 _24062_ (.A1_N(_13736_),
    .A2_N(_13742_),
    .B1(_13741_),
    .B2(_13744_),
    .Y(_14165_));
 sky130_fd_sc_hd__a2bb2o_1 _24063_ (.A1_N(_13736_),
    .A2_N(_13742_),
    .B1(_13741_),
    .B2(_13744_),
    .X(_14166_));
 sky130_fd_sc_hd__and3_2 _24064_ (.A(_14156_),
    .B(_09578_),
    .C(_14146_),
    .X(_14167_));
 sky130_fd_sc_hd__a21oi_4 _24065_ (.A1(_14161_),
    .A2(_14164_),
    .B1(_14165_),
    .Y(_14168_));
 sky130_fd_sc_hd__a31o_2 _24066_ (.A1(_14161_),
    .A2(_14164_),
    .A3(_14165_),
    .B1(_09578_),
    .X(_14169_));
 sky130_fd_sc_hd__nor2_1 _24067_ (.A(_14168_),
    .B(_14169_),
    .Y(_14170_));
 sky130_fd_sc_hd__o22ai_4 _24068_ (.A1(_09579_),
    .A2(_14160_),
    .B1(_14168_),
    .B2(_14169_),
    .Y(_14171_));
 sky130_fd_sc_hd__o22a_1 _24069_ (.A1(_09579_),
    .A2(_14160_),
    .B1(_14168_),
    .B2(_14169_),
    .X(_14172_));
 sky130_fd_sc_hd__o22a_1 _24070_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_14167_),
    .B2(_14170_),
    .X(_14174_));
 sky130_fd_sc_hd__o21ai_2 _24071_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_14171_),
    .Y(_14175_));
 sky130_fd_sc_hd__o21ai_1 _24072_ (.A1(_14168_),
    .A2(_14169_),
    .B1(_10015_),
    .Y(_14176_));
 sky130_fd_sc_hd__o221ai_2 _24073_ (.A1(_09579_),
    .A2(_14160_),
    .B1(_14168_),
    .B2(_14169_),
    .C1(_10015_),
    .Y(_14177_));
 sky130_fd_sc_hd__a31o_1 _24074_ (.A1(_08907_),
    .A2(_13749_),
    .A3(_13752_),
    .B1(_13754_),
    .X(_14178_));
 sky130_fd_sc_hd__a32o_1 _24075_ (.A1(_13753_),
    .A2(_08896_),
    .A3(_08874_),
    .B1(_13757_),
    .B2(_13755_),
    .X(_14179_));
 sky130_fd_sc_hd__o2111ai_1 _24076_ (.A1(_14167_),
    .A2(_14176_),
    .B1(_14178_),
    .C1(_14175_),
    .D1(_13758_),
    .Y(_14180_));
 sky130_fd_sc_hd__a22o_1 _24077_ (.A1(_14175_),
    .A2(_14177_),
    .B1(_14178_),
    .B2(_13758_),
    .X(_14181_));
 sky130_fd_sc_hd__o211ai_2 _24078_ (.A1(_10474_),
    .A2(net138),
    .B1(_14180_),
    .C1(_14181_),
    .Y(_14182_));
 sky130_fd_sc_hd__a21o_1 _24079_ (.A1(_14175_),
    .A2(_14177_),
    .B1(_14179_),
    .X(_14183_));
 sky130_fd_sc_hd__o21ai_2 _24080_ (.A1(_10025_),
    .A2(_14171_),
    .B1(_14179_),
    .Y(_14185_));
 sky130_fd_sc_hd__o221ai_4 _24081_ (.A1(_10474_),
    .A2(net138),
    .B1(_14174_),
    .B2(_14185_),
    .C1(_14183_),
    .Y(_14186_));
 sky130_fd_sc_hd__o31a_1 _24082_ (.A1(_10480_),
    .A2(_14167_),
    .A3(_14170_),
    .B1(_14182_),
    .X(_14187_));
 sky130_fd_sc_hd__o21ai_1 _24083_ (.A1(_07888_),
    .A2(_13761_),
    .B1(_13769_),
    .Y(_14188_));
 sky130_fd_sc_hd__o2111ai_4 _24084_ (.A1(_10480_),
    .A2(_14172_),
    .B1(_14186_),
    .C1(_08852_),
    .D1(_08830_),
    .Y(_14189_));
 sky130_fd_sc_hd__o211ai_2 _24085_ (.A1(_14171_),
    .A2(_10480_),
    .B1(_08918_),
    .C1(_14182_),
    .Y(_14190_));
 sky130_fd_sc_hd__a22o_1 _24086_ (.A1(_13762_),
    .A2(_13769_),
    .B1(_14189_),
    .B2(_14190_),
    .X(_14191_));
 sky130_fd_sc_hd__a41oi_1 _24087_ (.A1(_13762_),
    .A2(_13769_),
    .A3(_14189_),
    .A4(_14190_),
    .B1(_10953_),
    .Y(_14192_));
 sky130_fd_sc_hd__o2bb2a_1 _24088_ (.A1_N(_14191_),
    .A2_N(_14192_),
    .B1(_10954_),
    .B2(_14187_),
    .X(_14193_));
 sky130_fd_sc_hd__a2bb2o_1 _24089_ (.A1_N(_10954_),
    .A2_N(_14187_),
    .B1(_14191_),
    .B2(_14192_),
    .X(_14194_));
 sky130_fd_sc_hd__o21ai_1 _24090_ (.A1(_07800_),
    .A2(_07822_),
    .B1(_14193_),
    .Y(_14196_));
 sky130_fd_sc_hd__o21ai_1 _24091_ (.A1(net368),
    .A2(_07866_),
    .B1(_14194_),
    .Y(_14197_));
 sky130_fd_sc_hd__nand2_1 _24092_ (.A(_14196_),
    .B(_14197_),
    .Y(_14198_));
 sky130_fd_sc_hd__a21oi_1 _24093_ (.A1(_13772_),
    .A2(_13773_),
    .B1(_13774_),
    .Y(_14199_));
 sky130_fd_sc_hd__a21oi_1 _24094_ (.A1(_07888_),
    .A2(_14194_),
    .B1(_14199_),
    .Y(_14200_));
 sky130_fd_sc_hd__a221oi_1 _24095_ (.A1(_14198_),
    .A2(_14199_),
    .B1(_14200_),
    .B2(_14196_),
    .C1(_11464_),
    .Y(_14201_));
 sky130_fd_sc_hd__a31o_1 _24096_ (.A1(_11460_),
    .A2(_11462_),
    .A3(_14193_),
    .B1(_14201_),
    .X(_14202_));
 sky130_fd_sc_hd__and3_1 _24097_ (.A(_14202_),
    .B(_07022_),
    .C(net376),
    .X(_14203_));
 sky130_fd_sc_hd__a21oi_1 _24098_ (.A1(net376),
    .A2(_07022_),
    .B1(_14202_),
    .Y(_14204_));
 sky130_fd_sc_hd__o32ai_2 _24099_ (.A1(net394),
    .A2(_06267_),
    .A3(_13779_),
    .B1(_13781_),
    .B2(_13783_),
    .Y(_14205_));
 sky130_fd_sc_hd__o21ai_1 _24100_ (.A1(_14203_),
    .A2(_14204_),
    .B1(_14205_),
    .Y(_14207_));
 sky130_fd_sc_hd__a21oi_1 _24101_ (.A1(_14207_),
    .A2(_11943_),
    .B1(_14202_),
    .Y(_14208_));
 sky130_fd_sc_hd__xor2_1 _24102_ (.A(_13789_),
    .B(_14208_),
    .X(net94));
 sky130_fd_sc_hd__a2111oi_2 _24103_ (.A1(_11943_),
    .A2(_14207_),
    .B1(_13340_),
    .C1(_14202_),
    .D1(_13785_),
    .Y(_14209_));
 sky130_fd_sc_hd__o311a_1 _24104_ (.A1(_03399_),
    .A2(net24),
    .A3(_10962_),
    .B1(_13794_),
    .C1(_13800_),
    .X(_14210_));
 sky130_fd_sc_hd__a31o_1 _24105_ (.A1(_11471_),
    .A2(_13794_),
    .A3(_13800_),
    .B1(_08732_),
    .X(_14211_));
 sky130_fd_sc_hd__or4_1 _24106_ (.A(_08732_),
    .B(net351),
    .C(_09807_),
    .D(_14210_),
    .X(_14212_));
 sky130_fd_sc_hd__a311o_1 _24107_ (.A1(_11471_),
    .A2(_13794_),
    .A3(_13800_),
    .B1(_10970_),
    .C1(_08732_),
    .X(_14213_));
 sky130_fd_sc_hd__o21ai_1 _24108_ (.A1(_08732_),
    .A2(_14210_),
    .B1(_10970_),
    .Y(_14214_));
 sky130_fd_sc_hd__and2_1 _24109_ (.A(_14213_),
    .B(_14214_),
    .X(_14215_));
 sky130_fd_sc_hd__nand2_1 _24110_ (.A(_14213_),
    .B(_14214_),
    .Y(_14217_));
 sky130_fd_sc_hd__o21ai_2 _24111_ (.A1(_13809_),
    .A2(_13814_),
    .B1(_13807_),
    .Y(_14218_));
 sky130_fd_sc_hd__a21oi_1 _24112_ (.A1(_13807_),
    .A2(_13817_),
    .B1(_14217_),
    .Y(_14219_));
 sky130_fd_sc_hd__nand2_2 _24113_ (.A(_14218_),
    .B(_14215_),
    .Y(_14220_));
 sky130_fd_sc_hd__o211ai_1 _24114_ (.A1(_13809_),
    .A2(_13814_),
    .B1(_14217_),
    .C1(_13807_),
    .Y(_14221_));
 sky130_fd_sc_hd__o21ai_1 _24115_ (.A1(net351),
    .A2(_09807_),
    .B1(_14221_),
    .Y(_14222_));
 sky130_fd_sc_hd__o221ai_4 _24116_ (.A1(net351),
    .A2(_09807_),
    .B1(_14215_),
    .B2(_14218_),
    .C1(_14220_),
    .Y(_14223_));
 sky130_fd_sc_hd__o22ai_1 _24117_ (.A1(net335),
    .A2(_14211_),
    .B1(_14222_),
    .B2(_14219_),
    .Y(_14224_));
 sky130_fd_sc_hd__a21oi_2 _24118_ (.A1(_14212_),
    .A2(_14223_),
    .B1(net332),
    .Y(_14225_));
 sky130_fd_sc_hd__a2bb2oi_1 _24119_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_14212_),
    .B2(_14223_),
    .Y(_14226_));
 sky130_fd_sc_hd__o21ai_1 _24120_ (.A1(_10487_),
    .A2(net166),
    .B1(_14224_),
    .Y(_14228_));
 sky130_fd_sc_hd__o221a_1 _24121_ (.A1(net335),
    .A2(_14211_),
    .B1(_14222_),
    .B2(_14219_),
    .C1(net150),
    .X(_14229_));
 sky130_fd_sc_hd__o221ai_1 _24122_ (.A1(net335),
    .A2(_14211_),
    .B1(_14222_),
    .B2(_14219_),
    .C1(net150),
    .Y(_14230_));
 sky130_fd_sc_hd__nand2_1 _24123_ (.A(_14228_),
    .B(_14230_),
    .Y(_14231_));
 sky130_fd_sc_hd__a31oi_4 _24124_ (.A1(_13825_),
    .A2(_13830_),
    .A3(_13831_),
    .B1(_13823_),
    .Y(_14232_));
 sky130_fd_sc_hd__o21ai_2 _24125_ (.A1(_14226_),
    .A2(_14229_),
    .B1(_14232_),
    .Y(_14233_));
 sky130_fd_sc_hd__o221a_1 _24126_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_14232_),
    .B2(_14231_),
    .C1(_14233_),
    .X(_14234_));
 sky130_fd_sc_hd__o221ai_4 _24127_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_14232_),
    .B2(_14231_),
    .C1(_14233_),
    .Y(_14235_));
 sky130_fd_sc_hd__a21oi_1 _24128_ (.A1(_11079_),
    .A2(_14224_),
    .B1(_14234_),
    .Y(_14236_));
 sky130_fd_sc_hd__o21a_1 _24129_ (.A1(_14225_),
    .A2(_14234_),
    .B1(_12703_),
    .X(_14237_));
 sky130_fd_sc_hd__or3_1 _24130_ (.A(net329),
    .B(net327),
    .C(_14236_),
    .X(_14239_));
 sky130_fd_sc_hd__o22a_1 _24131_ (.A1(net170),
    .A2(net169),
    .B1(_14225_),
    .B2(_14234_),
    .X(_14240_));
 sky130_fd_sc_hd__o22ai_2 _24132_ (.A1(net170),
    .A2(net169),
    .B1(_14225_),
    .B2(_14234_),
    .Y(_14241_));
 sky130_fd_sc_hd__nand3b_4 _24133_ (.A_N(_14225_),
    .B(_14235_),
    .C(net153),
    .Y(_14242_));
 sky130_fd_sc_hd__and3_1 _24134_ (.A(_12970_),
    .B(_12518_),
    .C(_12968_),
    .X(_14243_));
 sky130_fd_sc_hd__nand3_1 _24135_ (.A(_13845_),
    .B(_14243_),
    .C(_13401_),
    .Y(_14244_));
 sky130_fd_sc_hd__o211ai_4 _24136_ (.A1(_13842_),
    .A2(_13844_),
    .B1(_13847_),
    .C1(_14244_),
    .Y(_14245_));
 sky130_fd_sc_hd__o2111a_1 _24137_ (.A1(_12522_),
    .A2(_12524_),
    .B1(_13398_),
    .C1(_13400_),
    .D1(_14243_),
    .X(_14246_));
 sky130_fd_sc_hd__nand3_4 _24138_ (.A(_14246_),
    .B(_13847_),
    .C(_13845_),
    .Y(_14247_));
 sky130_fd_sc_hd__a22oi_1 _24139_ (.A1(_14241_),
    .A2(_14242_),
    .B1(_14245_),
    .B2(_14247_),
    .Y(_14248_));
 sky130_fd_sc_hd__a22o_1 _24140_ (.A1(_14241_),
    .A2(_14242_),
    .B1(_14245_),
    .B2(_14247_),
    .X(_14250_));
 sky130_fd_sc_hd__nand4_2 _24141_ (.A(_14241_),
    .B(_14242_),
    .C(_14245_),
    .D(_14247_),
    .Y(_14251_));
 sky130_fd_sc_hd__o21ai_1 _24142_ (.A1(net329),
    .A2(net327),
    .B1(_14251_),
    .Y(_14252_));
 sky130_fd_sc_hd__nand3_1 _24143_ (.A(_14250_),
    .B(_14251_),
    .C(net311),
    .Y(_14253_));
 sky130_fd_sc_hd__o22ai_2 _24144_ (.A1(net311),
    .A2(_14236_),
    .B1(_14248_),
    .B2(_14252_),
    .Y(_14254_));
 sky130_fd_sc_hd__and3_2 _24145_ (.A(_00022_),
    .B(_00044_),
    .C(_14254_),
    .X(_14255_));
 sky130_fd_sc_hd__a211o_2 _24146_ (.A1(_14239_),
    .A2(_14253_),
    .B1(_00011_),
    .C1(net321),
    .X(_14256_));
 sky130_fd_sc_hd__a21oi_1 _24147_ (.A1(_13414_),
    .A2(_13852_),
    .B1(_13857_),
    .Y(_14257_));
 sky130_fd_sc_hd__a31o_1 _24148_ (.A1(_13414_),
    .A2(_13852_),
    .A3(_13856_),
    .B1(_13857_),
    .X(_14258_));
 sky130_fd_sc_hd__a31oi_2 _24149_ (.A1(_13414_),
    .A2(_13852_),
    .A3(_13856_),
    .B1(_13857_),
    .Y(_14259_));
 sky130_fd_sc_hd__a311oi_4 _24150_ (.A1(_14250_),
    .A2(_14251_),
    .A3(net311),
    .B1(_09595_),
    .C1(_14237_),
    .Y(_14261_));
 sky130_fd_sc_hd__nand3_2 _24151_ (.A(_14253_),
    .B(net172),
    .C(_14239_),
    .Y(_14262_));
 sky130_fd_sc_hd__a2bb2oi_1 _24152_ (.A1_N(_09588_),
    .A2_N(_09590_),
    .B1(_14239_),
    .B2(_14253_),
    .Y(_14263_));
 sky130_fd_sc_hd__o21ai_4 _24153_ (.A1(_09588_),
    .A2(_09590_),
    .B1(_14254_),
    .Y(_14264_));
 sky130_fd_sc_hd__nand3_4 _24154_ (.A(_14264_),
    .B(_14258_),
    .C(_14262_),
    .Y(_14265_));
 sky130_fd_sc_hd__o22ai_4 _24155_ (.A1(_13855_),
    .A2(_14257_),
    .B1(_14261_),
    .B2(_14263_),
    .Y(_14266_));
 sky130_fd_sc_hd__o211ai_4 _24156_ (.A1(_00011_),
    .A2(net323),
    .B1(_14265_),
    .C1(_14266_),
    .Y(_14267_));
 sky130_fd_sc_hd__a31oi_4 _24157_ (.A1(_14265_),
    .A2(_14266_),
    .A3(net307),
    .B1(_14255_),
    .Y(_14268_));
 sky130_fd_sc_hd__a31o_1 _24158_ (.A1(_14265_),
    .A2(_14266_),
    .A3(net307),
    .B1(_14255_),
    .X(_14269_));
 sky130_fd_sc_hd__a311oi_4 _24159_ (.A1(_14265_),
    .A2(_14266_),
    .A3(net307),
    .B1(net173),
    .C1(_14255_),
    .Y(_14270_));
 sky130_fd_sc_hd__o211ai_4 _24160_ (.A1(_09136_),
    .A2(_09138_),
    .B1(_14256_),
    .C1(_14267_),
    .Y(_14272_));
 sky130_fd_sc_hd__a2bb2oi_4 _24161_ (.A1_N(_09134_),
    .A2_N(_09135_),
    .B1(_14256_),
    .B2(_14267_),
    .Y(_14273_));
 sky130_fd_sc_hd__a2bb2o_1 _24162_ (.A1_N(_09134_),
    .A2_N(_09135_),
    .B1(_14256_),
    .B2(_14267_),
    .X(_14274_));
 sky130_fd_sc_hd__nor2_1 _24163_ (.A(_14270_),
    .B(_14273_),
    .Y(_14275_));
 sky130_fd_sc_hd__o211ai_4 _24164_ (.A1(net199),
    .A2(_13423_),
    .B1(_13870_),
    .C1(_13874_),
    .Y(_14276_));
 sky130_fd_sc_hd__o21ai_1 _24165_ (.A1(net175),
    .A2(_13868_),
    .B1(_14276_),
    .Y(_14277_));
 sky130_fd_sc_hd__nand4_1 _24166_ (.A(_13870_),
    .B(_13880_),
    .C(_14272_),
    .D(_14274_),
    .Y(_14278_));
 sky130_fd_sc_hd__o221ai_2 _24167_ (.A1(net175),
    .A2(_13868_),
    .B1(_14270_),
    .B2(_14273_),
    .C1(_14276_),
    .Y(_14279_));
 sky130_fd_sc_hd__nand3_2 _24168_ (.A(_14278_),
    .B(_14279_),
    .C(net278),
    .Y(_14280_));
 sky130_fd_sc_hd__o21ai_1 _24169_ (.A1(_14270_),
    .A2(_14273_),
    .B1(_14277_),
    .Y(_14281_));
 sky130_fd_sc_hd__o221ai_4 _24170_ (.A1(_13868_),
    .A2(net175),
    .B1(net174),
    .B2(_14268_),
    .C1(_14276_),
    .Y(_14283_));
 sky130_fd_sc_hd__o221ai_4 _24171_ (.A1(net304),
    .A2(_01951_),
    .B1(_14270_),
    .B2(_14283_),
    .C1(_14281_),
    .Y(_14284_));
 sky130_fd_sc_hd__o31a_2 _24172_ (.A1(net304),
    .A2(_01951_),
    .A3(_14268_),
    .B1(_14284_),
    .X(_14285_));
 sky130_fd_sc_hd__o211ai_4 _24173_ (.A1(_14269_),
    .A2(net278),
    .B1(net175),
    .C1(_14280_),
    .Y(_14286_));
 sky130_fd_sc_hd__o211ai_4 _24174_ (.A1(net278),
    .A2(_14268_),
    .B1(net177),
    .C1(_14284_),
    .Y(_14287_));
 sky130_fd_sc_hd__nand2_2 _24175_ (.A(_14286_),
    .B(_14287_),
    .Y(_14288_));
 sky130_fd_sc_hd__o2bb2ai_1 _24176_ (.A1_N(_13899_),
    .A2_N(_13902_),
    .B1(net199),
    .B2(_13884_),
    .Y(_14289_));
 sky130_fd_sc_hd__o21ai_1 _24177_ (.A1(net198),
    .A2(_13883_),
    .B1(_13902_),
    .Y(_14290_));
 sky130_fd_sc_hd__o22ai_1 _24178_ (.A1(net199),
    .A2(_13884_),
    .B1(_14290_),
    .B2(_13897_),
    .Y(_14291_));
 sky130_fd_sc_hd__a31oi_2 _24179_ (.A1(_13889_),
    .A2(_13899_),
    .A3(_13902_),
    .B1(_13885_),
    .Y(_14292_));
 sky130_fd_sc_hd__o2111ai_4 _24180_ (.A1(net198),
    .A2(_13883_),
    .B1(_14286_),
    .C1(_14287_),
    .D1(_14289_),
    .Y(_14294_));
 sky130_fd_sc_hd__o2bb2ai_2 _24181_ (.A1_N(_14286_),
    .A2_N(_14287_),
    .B1(_13897_),
    .B2(_13907_),
    .Y(_14295_));
 sky130_fd_sc_hd__o221ai_4 _24182_ (.A1(net199),
    .A2(_13884_),
    .B1(_13891_),
    .B2(_13904_),
    .C1(_14288_),
    .Y(_14296_));
 sky130_fd_sc_hd__o211a_2 _24183_ (.A1(_14269_),
    .A2(net278),
    .B1(_04040_),
    .C1(_14280_),
    .X(_14297_));
 sky130_fd_sc_hd__o221a_1 _24184_ (.A1(net302),
    .A2(_04019_),
    .B1(_13885_),
    .B2(_14295_),
    .C1(_14294_),
    .X(_14298_));
 sky130_fd_sc_hd__o221ai_4 _24185_ (.A1(net302),
    .A2(_04019_),
    .B1(_13885_),
    .B2(_14295_),
    .C1(_14294_),
    .Y(_14299_));
 sky130_fd_sc_hd__a31o_1 _24186_ (.A1(_14294_),
    .A2(_14296_),
    .A3(net277),
    .B1(_14297_),
    .X(_14300_));
 sky130_fd_sc_hd__a31oi_4 _24187_ (.A1(_14294_),
    .A2(_14296_),
    .A3(net277),
    .B1(_14297_),
    .Y(_14301_));
 sky130_fd_sc_hd__o22a_2 _24188_ (.A1(_05228_),
    .A2(_05230_),
    .B1(_14297_),
    .B2(_14298_),
    .X(_14302_));
 sky130_fd_sc_hd__or3_1 _24189_ (.A(net296),
    .B(_05232_),
    .C(_14301_),
    .X(_14303_));
 sky130_fd_sc_hd__and3_1 _24190_ (.A(_12581_),
    .B(_13038_),
    .C(_13039_),
    .X(_14305_));
 sky130_fd_sc_hd__nor3b_1 _24191_ (.A(_13469_),
    .B(_13472_),
    .C_N(_14305_),
    .Y(_14306_));
 sky130_fd_sc_hd__nand3_2 _24192_ (.A(_13917_),
    .B(_14305_),
    .C(_13474_),
    .Y(_14307_));
 sky130_fd_sc_hd__o211a_1 _24193_ (.A1(_13922_),
    .A2(_13916_),
    .B1(_13918_),
    .C1(_14307_),
    .X(_14308_));
 sky130_fd_sc_hd__o211ai_4 _24194_ (.A1(_13922_),
    .A2(_13916_),
    .B1(_13918_),
    .C1(_14307_),
    .Y(_14309_));
 sky130_fd_sc_hd__nand4_4 _24195_ (.A(_14306_),
    .B(_13918_),
    .C(_13917_),
    .D(_12592_),
    .Y(_14310_));
 sky130_fd_sc_hd__a41o_1 _24196_ (.A1(_12592_),
    .A2(_13917_),
    .A3(_13918_),
    .A4(_14306_),
    .B1(_14308_),
    .X(_14311_));
 sky130_fd_sc_hd__a21oi_2 _24197_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_14301_),
    .Y(_14312_));
 sky130_fd_sc_hd__o22ai_4 _24198_ (.A1(_08307_),
    .A2(net216),
    .B1(_14297_),
    .B2(_14298_),
    .Y(_14313_));
 sky130_fd_sc_hd__o221a_1 _24199_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_14285_),
    .B2(_04029_),
    .C1(_14299_),
    .X(_14314_));
 sky130_fd_sc_hd__o221ai_4 _24200_ (.A1(_08311_),
    .A2(_08312_),
    .B1(_14285_),
    .B2(_04029_),
    .C1(_14299_),
    .Y(_14316_));
 sky130_fd_sc_hd__a22oi_1 _24201_ (.A1(_14309_),
    .A2(_14310_),
    .B1(_14313_),
    .B2(_14316_),
    .Y(_14317_));
 sky130_fd_sc_hd__o2bb2ai_4 _24202_ (.A1_N(_14309_),
    .A2_N(_14310_),
    .B1(_14312_),
    .B2(_14314_),
    .Y(_14318_));
 sky130_fd_sc_hd__and4_1 _24203_ (.A(_14309_),
    .B(_14310_),
    .C(_14313_),
    .D(_14316_),
    .X(_14319_));
 sky130_fd_sc_hd__nand4_4 _24204_ (.A(_14309_),
    .B(_14310_),
    .C(_14313_),
    .D(_14316_),
    .Y(_14320_));
 sky130_fd_sc_hd__nand3_1 _24205_ (.A(_14318_),
    .B(_14320_),
    .C(net271),
    .Y(_14321_));
 sky130_fd_sc_hd__o22ai_2 _24206_ (.A1(net296),
    .A2(_05232_),
    .B1(_14317_),
    .B2(_14319_),
    .Y(_14322_));
 sky130_fd_sc_hd__a31oi_4 _24207_ (.A1(_14318_),
    .A2(_14320_),
    .A3(net271),
    .B1(_14302_),
    .Y(_14323_));
 sky130_fd_sc_hd__o221a_2 _24208_ (.A1(_05478_),
    .A2(_05479_),
    .B1(_14300_),
    .B2(net271),
    .C1(_14322_),
    .X(_14324_));
 sky130_fd_sc_hd__or3_4 _24209_ (.A(net270),
    .B(net268),
    .C(_14323_),
    .X(_14325_));
 sky130_fd_sc_hd__a31o_1 _24210_ (.A1(_14318_),
    .A2(_14320_),
    .A3(net271),
    .B1(_07936_),
    .X(_14327_));
 sky130_fd_sc_hd__a311oi_4 _24211_ (.A1(_14318_),
    .A2(_14320_),
    .A3(net271),
    .B1(_07936_),
    .C1(_14302_),
    .Y(_14328_));
 sky130_fd_sc_hd__nand3_1 _24212_ (.A(_14321_),
    .B(_07935_),
    .C(_14303_),
    .Y(_14329_));
 sky130_fd_sc_hd__a2bb2oi_2 _24213_ (.A1_N(_07928_),
    .A2_N(_07930_),
    .B1(_14303_),
    .B2(_14321_),
    .Y(_14330_));
 sky130_fd_sc_hd__o221ai_4 _24214_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_14300_),
    .B2(net271),
    .C1(_14322_),
    .Y(_14331_));
 sky130_fd_sc_hd__a31o_1 _24215_ (.A1(_13488_),
    .A2(_13929_),
    .A3(_13933_),
    .B1(_13934_),
    .X(_14332_));
 sky130_fd_sc_hd__a31oi_4 _24216_ (.A1(_13488_),
    .A2(_13929_),
    .A3(_13933_),
    .B1(_13934_),
    .Y(_14333_));
 sky130_fd_sc_hd__o21ai_4 _24217_ (.A1(_14328_),
    .A2(_14330_),
    .B1(_14333_),
    .Y(_14334_));
 sky130_fd_sc_hd__o211ai_4 _24218_ (.A1(_14302_),
    .A2(_14327_),
    .B1(_14332_),
    .C1(_14331_),
    .Y(_14335_));
 sky130_fd_sc_hd__o311a_1 _24219_ (.A1(_14328_),
    .A2(_14330_),
    .A3(_14333_),
    .B1(net245),
    .C1(_14334_),
    .X(_14336_));
 sky130_fd_sc_hd__nand3_2 _24220_ (.A(_14334_),
    .B(_14335_),
    .C(net245),
    .Y(_14338_));
 sky130_fd_sc_hd__a31o_2 _24221_ (.A1(_14334_),
    .A2(_14335_),
    .A3(net245),
    .B1(_14324_),
    .X(_14339_));
 sky130_fd_sc_hd__o221ai_4 _24222_ (.A1(net227),
    .A2(_13501_),
    .B1(_07246_),
    .B2(_13945_),
    .C1(_13951_),
    .Y(_14340_));
 sky130_fd_sc_hd__a22o_1 _24223_ (.A1(_07246_),
    .A2(_13945_),
    .B1(_13951_),
    .B2(_13505_),
    .X(_14341_));
 sky130_fd_sc_hd__a31oi_2 _24224_ (.A1(_14334_),
    .A2(_14335_),
    .A3(net245),
    .B1(net202),
    .Y(_14342_));
 sky130_fd_sc_hd__a311oi_4 _24225_ (.A1(_14334_),
    .A2(_14335_),
    .A3(net245),
    .B1(net202),
    .C1(_14324_),
    .Y(_14343_));
 sky130_fd_sc_hd__o211ai_4 _24226_ (.A1(net245),
    .A2(_14323_),
    .B1(_07564_),
    .C1(_14338_),
    .Y(_14344_));
 sky130_fd_sc_hd__a2bb2oi_4 _24227_ (.A1_N(net221),
    .A2_N(net220),
    .B1(_14325_),
    .B2(_14338_),
    .Y(_14345_));
 sky130_fd_sc_hd__o22ai_2 _24228_ (.A1(net221),
    .A2(net220),
    .B1(_14324_),
    .B2(_14336_),
    .Y(_14346_));
 sky130_fd_sc_hd__a21oi_1 _24229_ (.A1(_14325_),
    .A2(_14342_),
    .B1(_14345_),
    .Y(_14347_));
 sky130_fd_sc_hd__o2111ai_4 _24230_ (.A1(_13945_),
    .A2(_07246_),
    .B1(_14344_),
    .C1(_14341_),
    .D1(_14346_),
    .Y(_14349_));
 sky130_fd_sc_hd__o2bb2ai_1 _24231_ (.A1_N(_13947_),
    .A2_N(_14341_),
    .B1(_14343_),
    .B2(_14345_),
    .Y(_14350_));
 sky130_fd_sc_hd__o211ai_4 _24232_ (.A1(_05750_),
    .A2(net264),
    .B1(_14349_),
    .C1(_14350_),
    .Y(_14351_));
 sky130_fd_sc_hd__a211o_1 _24233_ (.A1(_14325_),
    .A2(_14338_),
    .B1(net265),
    .C1(net264),
    .X(_14352_));
 sky130_fd_sc_hd__o2111ai_1 _24234_ (.A1(net223),
    .A2(_13944_),
    .B1(_14340_),
    .C1(_14344_),
    .D1(_14346_),
    .Y(_14353_));
 sky130_fd_sc_hd__o2bb2ai_1 _24235_ (.A1_N(_13948_),
    .A2_N(_14340_),
    .B1(_14343_),
    .B2(_14345_),
    .Y(_14354_));
 sky130_fd_sc_hd__nand3_2 _24236_ (.A(_14353_),
    .B(_14354_),
    .C(net243),
    .Y(_14355_));
 sky130_fd_sc_hd__o31a_1 _24237_ (.A1(net243),
    .A2(_14324_),
    .A3(_14336_),
    .B1(_14351_),
    .X(_14356_));
 sky130_fd_sc_hd__o21ai_4 _24238_ (.A1(net243),
    .A2(_14339_),
    .B1(_14351_),
    .Y(_14357_));
 sky130_fd_sc_hd__a2bb2oi_1 _24239_ (.A1_N(_07242_),
    .A2_N(net248),
    .B1(_14352_),
    .B2(_14355_),
    .Y(_14358_));
 sky130_fd_sc_hd__o211ai_4 _24240_ (.A1(_14339_),
    .A2(net243),
    .B1(net222),
    .C1(_14351_),
    .Y(_14360_));
 sky130_fd_sc_hd__o211a_1 _24241_ (.A1(_07244_),
    .A2(net247),
    .B1(_14352_),
    .C1(_14355_),
    .X(_14361_));
 sky130_fd_sc_hd__nand3_4 _24242_ (.A(_14355_),
    .B(_07246_),
    .C(_14352_),
    .Y(_14362_));
 sky130_fd_sc_hd__nand2_1 _24243_ (.A(_14360_),
    .B(_14362_),
    .Y(_14363_));
 sky130_fd_sc_hd__o2bb2ai_2 _24244_ (.A1_N(_13968_),
    .A2_N(_13969_),
    .B1(net227),
    .B2(_13960_),
    .Y(_14364_));
 sky130_fd_sc_hd__nand3_2 _24245_ (.A(_13968_),
    .B(_13969_),
    .C(_13977_),
    .Y(_14365_));
 sky130_fd_sc_hd__a31oi_4 _24246_ (.A1(_13968_),
    .A2(_13969_),
    .A3(_13977_),
    .B1(_13972_),
    .Y(_14366_));
 sky130_fd_sc_hd__a22oi_4 _24247_ (.A1(_14360_),
    .A2(_14362_),
    .B1(_14364_),
    .B2(_13977_),
    .Y(_14367_));
 sky130_fd_sc_hd__o21ai_2 _24248_ (.A1(_14358_),
    .A2(_14361_),
    .B1(_14366_),
    .Y(_14368_));
 sky130_fd_sc_hd__o2111ai_4 _24249_ (.A1(_06924_),
    .A2(_13961_),
    .B1(_14360_),
    .C1(_14362_),
    .D1(_14364_),
    .Y(_14369_));
 sky130_fd_sc_hd__o22ai_4 _24250_ (.A1(net260),
    .A2(net258),
    .B1(_14363_),
    .B2(_14366_),
    .Y(_14371_));
 sky130_fd_sc_hd__o211ai_2 _24251_ (.A1(net260),
    .A2(net258),
    .B1(_14368_),
    .C1(_14369_),
    .Y(_14372_));
 sky130_fd_sc_hd__or3_4 _24252_ (.A(net260),
    .B(net258),
    .C(_14357_),
    .X(_14373_));
 sky130_fd_sc_hd__o22ai_4 _24253_ (.A1(net240),
    .A2(_14357_),
    .B1(_14367_),
    .B2(_14371_),
    .Y(_14374_));
 sky130_fd_sc_hd__inv_2 _24254_ (.A(_14374_),
    .Y(_14375_));
 sky130_fd_sc_hd__a22oi_4 _24255_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_14372_),
    .B2(_14373_),
    .Y(_14376_));
 sky130_fd_sc_hd__o21ai_2 _24256_ (.A1(_06914_),
    .A2(net250),
    .B1(_14374_),
    .Y(_14377_));
 sky130_fd_sc_hd__a31oi_4 _24257_ (.A1(net240),
    .A2(_14368_),
    .A3(_14369_),
    .B1(_06924_),
    .Y(_14378_));
 sky130_fd_sc_hd__o221ai_4 _24258_ (.A1(net240),
    .A2(_14357_),
    .B1(_14367_),
    .B2(_14371_),
    .C1(net227),
    .Y(_14379_));
 sky130_fd_sc_hd__a21oi_1 _24259_ (.A1(_14373_),
    .A2(_14378_),
    .B1(_14376_),
    .Y(_14380_));
 sky130_fd_sc_hd__and3_1 _24260_ (.A(_13129_),
    .B(_12656_),
    .C(_13127_),
    .X(_14382_));
 sky130_fd_sc_hd__nand3_1 _24261_ (.A(_13991_),
    .B(_14382_),
    .C(_13557_),
    .Y(_14383_));
 sky130_fd_sc_hd__o211ai_4 _24262_ (.A1(_13995_),
    .A2(_13990_),
    .B1(_13993_),
    .C1(_14383_),
    .Y(_14384_));
 sky130_fd_sc_hd__and4_1 _24263_ (.A(_14382_),
    .B(_13556_),
    .C(_13554_),
    .D(_12664_),
    .X(_14385_));
 sky130_fd_sc_hd__nand3_4 _24264_ (.A(_14385_),
    .B(_13993_),
    .C(_13991_),
    .Y(_14386_));
 sky130_fd_sc_hd__nand2_2 _24265_ (.A(_14384_),
    .B(_14386_),
    .Y(_14387_));
 sky130_fd_sc_hd__a221oi_4 _24266_ (.A1(_14373_),
    .A2(_14378_),
    .B1(_14384_),
    .B2(_14386_),
    .C1(_14376_),
    .Y(_14388_));
 sky130_fd_sc_hd__o22ai_2 _24267_ (.A1(net239),
    .A2(_06292_),
    .B1(_14380_),
    .B2(_14387_),
    .Y(_14389_));
 sky130_fd_sc_hd__a22o_1 _24268_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_14372_),
    .B2(_14373_),
    .X(_14390_));
 sky130_fd_sc_hd__inv_2 _24269_ (.A(_14390_),
    .Y(_14391_));
 sky130_fd_sc_hd__a22o_1 _24270_ (.A1(_14377_),
    .A2(_14379_),
    .B1(_14384_),
    .B2(_14386_),
    .X(_14393_));
 sky130_fd_sc_hd__nand3_2 _24271_ (.A(_14379_),
    .B(_14384_),
    .C(_14386_),
    .Y(_14394_));
 sky130_fd_sc_hd__o2111ai_4 _24272_ (.A1(_06924_),
    .A2(_14374_),
    .B1(_14377_),
    .C1(_14384_),
    .D1(_14386_),
    .Y(_14395_));
 sky130_fd_sc_hd__nand3_2 _24273_ (.A(_14393_),
    .B(_14395_),
    .C(net214),
    .Y(_14396_));
 sky130_fd_sc_hd__o221a_2 _24274_ (.A1(net214),
    .A2(_14374_),
    .B1(_14388_),
    .B2(_14389_),
    .C1(_06613_),
    .X(_14397_));
 sky130_fd_sc_hd__a211o_2 _24275_ (.A1(_14390_),
    .A2(_14396_),
    .B1(net238),
    .C1(_06610_),
    .X(_14398_));
 sky130_fd_sc_hd__a311oi_2 _24276_ (.A1(_14393_),
    .A2(_14395_),
    .A3(net214),
    .B1(net233),
    .C1(_14391_),
    .Y(_14399_));
 sky130_fd_sc_hd__nand3_4 _24277_ (.A(_14396_),
    .B(net235),
    .C(_14390_),
    .Y(_14400_));
 sky130_fd_sc_hd__o221ai_4 _24278_ (.A1(net214),
    .A2(_14374_),
    .B1(_14388_),
    .B2(_14389_),
    .C1(net233),
    .Y(_14401_));
 sky130_fd_sc_hd__o22a_1 _24279_ (.A1(_06314_),
    .A2(_14003_),
    .B1(_14005_),
    .B2(_13567_),
    .X(_14402_));
 sky130_fd_sc_hd__o32a_1 _24280_ (.A1(net284),
    .A2(net282),
    .A3(_14004_),
    .B1(_14007_),
    .B2(_14011_),
    .X(_14404_));
 sky130_fd_sc_hd__a21oi_1 _24281_ (.A1(_14007_),
    .A2(_14010_),
    .B1(_14011_),
    .Y(_14405_));
 sky130_fd_sc_hd__o2bb2ai_4 _24282_ (.A1_N(_14400_),
    .A2_N(_14401_),
    .B1(_14402_),
    .B2(_14009_),
    .Y(_14406_));
 sky130_fd_sc_hd__nand3_4 _24283_ (.A(_14404_),
    .B(_14401_),
    .C(_14400_),
    .Y(_14407_));
 sky130_fd_sc_hd__and3_1 _24284_ (.A(_14406_),
    .B(_14407_),
    .C(net210),
    .X(_14408_));
 sky130_fd_sc_hd__nand3_2 _24285_ (.A(_14406_),
    .B(_14407_),
    .C(net210),
    .Y(_14409_));
 sky130_fd_sc_hd__a31o_2 _24286_ (.A1(_14406_),
    .A2(_14407_),
    .A3(net210),
    .B1(_14397_),
    .X(_14410_));
 sky130_fd_sc_hd__and3_1 _24287_ (.A(_06904_),
    .B(_14398_),
    .C(_14409_),
    .X(_14411_));
 sky130_fd_sc_hd__o311a_1 _24288_ (.A1(_05765_),
    .A2(_05766_),
    .A3(_13583_),
    .B1(_13609_),
    .C1(_14024_),
    .X(_14412_));
 sky130_fd_sc_hd__a2bb2oi_2 _24289_ (.A1_N(_06014_),
    .A2_N(_14022_),
    .B1(_13609_),
    .B2(_13586_),
    .Y(_14413_));
 sky130_fd_sc_hd__a31oi_2 _24290_ (.A1(_13586_),
    .A2(_13609_),
    .A3(_14024_),
    .B1(_14025_),
    .Y(_14415_));
 sky130_fd_sc_hd__a31oi_1 _24291_ (.A1(_14406_),
    .A2(_14407_),
    .A3(net210),
    .B1(net252),
    .Y(_14416_));
 sky130_fd_sc_hd__a311oi_4 _24292_ (.A1(_14406_),
    .A2(_14407_),
    .A3(net210),
    .B1(_14397_),
    .C1(net252),
    .Y(_14417_));
 sky130_fd_sc_hd__a311o_2 _24293_ (.A1(_14406_),
    .A2(_14407_),
    .A3(net210),
    .B1(_14397_),
    .C1(net252),
    .X(_14418_));
 sky130_fd_sc_hd__a2bb2oi_4 _24294_ (.A1_N(net284),
    .A2_N(net282),
    .B1(_14398_),
    .B2(_14409_),
    .Y(_14419_));
 sky130_fd_sc_hd__o21ai_2 _24295_ (.A1(net284),
    .A2(net282),
    .B1(_14410_),
    .Y(_14420_));
 sky130_fd_sc_hd__o211ai_4 _24296_ (.A1(_14025_),
    .A2(_14412_),
    .B1(_14418_),
    .C1(_14420_),
    .Y(_14421_));
 sky130_fd_sc_hd__o22ai_4 _24297_ (.A1(_14023_),
    .A2(_14413_),
    .B1(_14417_),
    .B2(_14419_),
    .Y(_14422_));
 sky130_fd_sc_hd__o211ai_2 _24298_ (.A1(net231),
    .A2(net228),
    .B1(_14421_),
    .C1(_14422_),
    .Y(_14423_));
 sky130_fd_sc_hd__a211o_1 _24299_ (.A1(_14398_),
    .A2(_14409_),
    .B1(net231),
    .C1(net228),
    .X(_14424_));
 sky130_fd_sc_hd__o211ai_1 _24300_ (.A1(_14023_),
    .A2(_14413_),
    .B1(_14418_),
    .C1(_14420_),
    .Y(_14426_));
 sky130_fd_sc_hd__o22ai_1 _24301_ (.A1(_14025_),
    .A2(_14412_),
    .B1(_14417_),
    .B2(_14419_),
    .Y(_14427_));
 sky130_fd_sc_hd__nand3_2 _24302_ (.A(_14426_),
    .B(_14427_),
    .C(net208),
    .Y(_14428_));
 sky130_fd_sc_hd__a31o_2 _24303_ (.A1(_14421_),
    .A2(_14422_),
    .A3(net208),
    .B1(_14411_),
    .X(_14429_));
 sky130_fd_sc_hd__inv_2 _24304_ (.A(_14429_),
    .Y(_14430_));
 sky130_fd_sc_hd__nand2_1 _24305_ (.A(_14429_),
    .B(_07232_),
    .Y(_14431_));
 sky130_fd_sc_hd__a311oi_4 _24306_ (.A1(_14421_),
    .A2(_14422_),
    .A3(net208),
    .B1(_14411_),
    .C1(net254),
    .Y(_14432_));
 sky130_fd_sc_hd__o211ai_4 _24307_ (.A1(_14410_),
    .A2(net208),
    .B1(_06014_),
    .C1(_14423_),
    .Y(_14433_));
 sky130_fd_sc_hd__o211a_2 _24308_ (.A1(_06011_),
    .A2(_06012_),
    .B1(_14424_),
    .C1(_14428_),
    .X(_14434_));
 sky130_fd_sc_hd__o211ai_4 _24309_ (.A1(net285),
    .A2(_06012_),
    .B1(_14424_),
    .C1(_14428_),
    .Y(_14435_));
 sky130_fd_sc_hd__nand2_1 _24310_ (.A(_14433_),
    .B(_14435_),
    .Y(_14437_));
 sky130_fd_sc_hd__a22o_1 _24311_ (.A1(_05768_),
    .A2(_14037_),
    .B1(_14046_),
    .B2(_14047_),
    .X(_14438_));
 sky130_fd_sc_hd__a31oi_2 _24312_ (.A1(_14040_),
    .A2(_14046_),
    .A3(_14047_),
    .B1(_14038_),
    .Y(_14439_));
 sky130_fd_sc_hd__nand4_2 _24313_ (.A(_14039_),
    .B(_14055_),
    .C(_14433_),
    .D(_14435_),
    .Y(_14440_));
 sky130_fd_sc_hd__o2bb2ai_1 _24314_ (.A1_N(_14039_),
    .A2_N(_14055_),
    .B1(_14432_),
    .B2(_14434_),
    .Y(_14441_));
 sky130_fd_sc_hd__o211ai_4 _24315_ (.A1(net207),
    .A2(net206),
    .B1(_14440_),
    .C1(_14441_),
    .Y(_14442_));
 sky130_fd_sc_hd__o311a_1 _24316_ (.A1(net208),
    .A2(_14397_),
    .A3(_14408_),
    .B1(_07232_),
    .C1(_14423_),
    .X(_14443_));
 sky130_fd_sc_hd__a22oi_4 _24317_ (.A1(_14433_),
    .A2(_14435_),
    .B1(_14438_),
    .B2(_14040_),
    .Y(_14444_));
 sky130_fd_sc_hd__o22ai_4 _24318_ (.A1(net207),
    .A2(net206),
    .B1(_14437_),
    .B2(_14439_),
    .Y(_14445_));
 sky130_fd_sc_hd__o22ai_4 _24319_ (.A1(_07233_),
    .A2(_14429_),
    .B1(_14444_),
    .B2(_14445_),
    .Y(_14446_));
 sky130_fd_sc_hd__inv_2 _24320_ (.A(_14446_),
    .Y(_14448_));
 sky130_fd_sc_hd__o211a_1 _24321_ (.A1(_14430_),
    .A2(_07233_),
    .B1(_05768_),
    .C1(_14442_),
    .X(_14449_));
 sky130_fd_sc_hd__o211ai_4 _24322_ (.A1(_14430_),
    .A2(_07233_),
    .B1(_05768_),
    .C1(_14442_),
    .Y(_14450_));
 sky130_fd_sc_hd__o21ai_1 _24323_ (.A1(_14444_),
    .A2(_14445_),
    .B1(net263),
    .Y(_14451_));
 sky130_fd_sc_hd__o221a_2 _24324_ (.A1(_07233_),
    .A2(_14429_),
    .B1(_14444_),
    .B2(_14445_),
    .C1(net263),
    .X(_14452_));
 sky130_fd_sc_hd__a21o_1 _24325_ (.A1(_14431_),
    .A2(_14442_),
    .B1(_05768_),
    .X(_14453_));
 sky130_fd_sc_hd__o21ai_2 _24326_ (.A1(_14443_),
    .A2(_14451_),
    .B1(_14450_),
    .Y(_14454_));
 sky130_fd_sc_hd__nand4_2 _24327_ (.A(_12721_),
    .B(_12723_),
    .C(_13201_),
    .D(_13203_),
    .Y(_14455_));
 sky130_fd_sc_hd__a211oi_4 _24328_ (.A1(_13615_),
    .A2(_13637_),
    .B1(_14455_),
    .C1(_13640_),
    .Y(_14456_));
 sky130_fd_sc_hd__nand2_1 _24329_ (.A(_14062_),
    .B(_14456_),
    .Y(_14457_));
 sky130_fd_sc_hd__o211a_1 _24330_ (.A1(_14067_),
    .A2(_14061_),
    .B1(_14064_),
    .C1(_14457_),
    .X(_14459_));
 sky130_fd_sc_hd__o211ai_4 _24331_ (.A1(_14067_),
    .A2(_14061_),
    .B1(_14064_),
    .C1(_14457_),
    .Y(_14460_));
 sky130_fd_sc_hd__nand3_1 _24332_ (.A(_14062_),
    .B(_14456_),
    .C(_14064_),
    .Y(_14461_));
 sky130_fd_sc_hd__nand4_4 _24333_ (.A(_14062_),
    .B(_14456_),
    .C(_14064_),
    .D(_12730_),
    .Y(_14462_));
 sky130_fd_sc_hd__a41o_1 _24334_ (.A1(_12730_),
    .A2(_14062_),
    .A3(_14064_),
    .A4(_14456_),
    .B1(_14459_),
    .X(_14463_));
 sky130_fd_sc_hd__a21oi_4 _24335_ (.A1(_14460_),
    .A2(_14462_),
    .B1(_14454_),
    .Y(_14464_));
 sky130_fd_sc_hd__o221ai_4 _24336_ (.A1(_14461_),
    .A2(_12731_),
    .B1(_14449_),
    .B2(_14452_),
    .C1(_14460_),
    .Y(_14465_));
 sky130_fd_sc_hd__o21ai_4 _24337_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_14465_),
    .Y(_14466_));
 sky130_fd_sc_hd__and3_1 _24338_ (.A(_07550_),
    .B(_14431_),
    .C(_14442_),
    .X(_14467_));
 sky130_fd_sc_hd__or3b_1 _24339_ (.A(_07544_),
    .B(_07546_),
    .C_N(_14446_),
    .X(_14468_));
 sky130_fd_sc_hd__a22o_1 _24340_ (.A1(_14450_),
    .A2(_14453_),
    .B1(_14460_),
    .B2(_14462_),
    .X(_00001_));
 sky130_fd_sc_hd__o21ai_1 _24341_ (.A1(_05768_),
    .A2(_14446_),
    .B1(_14462_),
    .Y(_00002_));
 sky130_fd_sc_hd__o211ai_1 _24342_ (.A1(_14446_),
    .A2(_05768_),
    .B1(_14462_),
    .C1(_14460_),
    .Y(_00003_));
 sky130_fd_sc_hd__o2111ai_2 _24343_ (.A1(_05768_),
    .A2(_14446_),
    .B1(_14450_),
    .C1(_14460_),
    .D1(_14462_),
    .Y(_00004_));
 sky130_fd_sc_hd__nand3_1 _24344_ (.A(_00001_),
    .B(_00004_),
    .C(net163),
    .Y(_00005_));
 sky130_fd_sc_hd__a31o_1 _24345_ (.A1(_00001_),
    .A2(_00004_),
    .A3(net163),
    .B1(_14467_),
    .X(_00006_));
 sky130_fd_sc_hd__o22ai_4 _24346_ (.A1(net163),
    .A2(_14446_),
    .B1(_14464_),
    .B2(_14466_),
    .Y(_00007_));
 sky130_fd_sc_hd__o221a_1 _24347_ (.A1(net163),
    .A2(_14446_),
    .B1(_14464_),
    .B2(_14466_),
    .C1(_07917_),
    .X(_00008_));
 sky130_fd_sc_hd__or3_2 _24348_ (.A(net183),
    .B(net182),
    .C(_00007_),
    .X(_00009_));
 sky130_fd_sc_hd__a31o_1 _24349_ (.A1(_00001_),
    .A2(_00004_),
    .A3(net163),
    .B1(net292),
    .X(_00010_));
 sky130_fd_sc_hd__nand3_4 _24350_ (.A(_00005_),
    .B(_05507_),
    .C(_14468_),
    .Y(_00012_));
 sky130_fd_sc_hd__o221ai_4 _24351_ (.A1(net163),
    .A2(_14446_),
    .B1(_14464_),
    .B2(_14466_),
    .C1(net292),
    .Y(_00013_));
 sky130_fd_sc_hd__o221a_1 _24352_ (.A1(_13650_),
    .A2(_04227_),
    .B1(net295),
    .B2(_14076_),
    .C1(_14080_),
    .X(_00014_));
 sky130_fd_sc_hd__o22a_1 _24353_ (.A1(_13651_),
    .A2(_14079_),
    .B1(_14077_),
    .B2(net294),
    .X(_00015_));
 sky130_fd_sc_hd__a21o_1 _24354_ (.A1(_14081_),
    .A2(_14083_),
    .B1(_14084_),
    .X(_00016_));
 sky130_fd_sc_hd__o31a_1 _24355_ (.A1(_13653_),
    .A2(_14078_),
    .A3(_14082_),
    .B1(_14086_),
    .X(_00017_));
 sky130_fd_sc_hd__a21oi_4 _24356_ (.A1(_00012_),
    .A2(_00013_),
    .B1(_00016_),
    .Y(_00018_));
 sky130_fd_sc_hd__o2bb2ai_2 _24357_ (.A1_N(_00012_),
    .A2_N(_00013_),
    .B1(_00014_),
    .B2(_14082_),
    .Y(_00019_));
 sky130_fd_sc_hd__o211a_1 _24358_ (.A1(_14084_),
    .A2(_00015_),
    .B1(_00013_),
    .C1(_00012_),
    .X(_00020_));
 sky130_fd_sc_hd__o211ai_4 _24359_ (.A1(_14084_),
    .A2(_00015_),
    .B1(_00013_),
    .C1(_00012_),
    .Y(_00021_));
 sky130_fd_sc_hd__a31o_1 _24360_ (.A1(_00012_),
    .A2(_00013_),
    .A3(_00016_),
    .B1(_07917_),
    .X(_00023_));
 sky130_fd_sc_hd__nand3_1 _24361_ (.A(_00019_),
    .B(_00021_),
    .C(net161),
    .Y(_00024_));
 sky130_fd_sc_hd__o22ai_2 _24362_ (.A1(net183),
    .A2(net182),
    .B1(_00018_),
    .B2(_00020_),
    .Y(_00025_));
 sky130_fd_sc_hd__o22ai_4 _24363_ (.A1(net161),
    .A2(_00007_),
    .B1(_00018_),
    .B2(_00023_),
    .Y(_00026_));
 sky130_fd_sc_hd__a311o_1 _24364_ (.A1(_00019_),
    .A2(_00021_),
    .A3(net161),
    .B1(net159),
    .C1(_00008_),
    .X(_00027_));
 sky130_fd_sc_hd__o221a_1 _24365_ (.A1(_13666_),
    .A2(_13678_),
    .B1(_04227_),
    .B2(_14094_),
    .C1(_13665_),
    .X(_00028_));
 sky130_fd_sc_hd__a21oi_1 _24366_ (.A1(_04227_),
    .A2(_14094_),
    .B1(_14102_),
    .Y(_00029_));
 sky130_fd_sc_hd__o21ai_2 _24367_ (.A1(_14102_),
    .A2(_14098_),
    .B1(_14097_),
    .Y(_00030_));
 sky130_fd_sc_hd__a32o_1 _24368_ (.A1(_04173_),
    .A2(_04195_),
    .A3(_14094_),
    .B1(_14097_),
    .B2(_14102_),
    .X(_00031_));
 sky130_fd_sc_hd__a311oi_4 _24369_ (.A1(_00019_),
    .A2(_00021_),
    .A3(net161),
    .B1(_00008_),
    .C1(net294),
    .Y(_00032_));
 sky130_fd_sc_hd__o221ai_4 _24370_ (.A1(net161),
    .A2(_00007_),
    .B1(_00018_),
    .B2(_00023_),
    .C1(net295),
    .Y(_00034_));
 sky130_fd_sc_hd__a2bb2oi_4 _24371_ (.A1_N(net318),
    .A2_N(net316),
    .B1(_00009_),
    .B2(_00024_),
    .Y(_00035_));
 sky130_fd_sc_hd__o221ai_4 _24372_ (.A1(net318),
    .A2(net315),
    .B1(net161),
    .B2(_00006_),
    .C1(_00025_),
    .Y(_00036_));
 sky130_fd_sc_hd__o211ai_2 _24373_ (.A1(_14098_),
    .A2(_00028_),
    .B1(_00034_),
    .C1(_00036_),
    .Y(_00037_));
 sky130_fd_sc_hd__o22ai_2 _24374_ (.A1(_14095_),
    .A2(_00029_),
    .B1(_00032_),
    .B2(_00035_),
    .Y(_00038_));
 sky130_fd_sc_hd__o211ai_4 _24375_ (.A1(_08296_),
    .A2(_08298_),
    .B1(_00037_),
    .C1(_00038_),
    .Y(_00039_));
 sky130_fd_sc_hd__o221a_1 _24376_ (.A1(_08293_),
    .A2(_08295_),
    .B1(_00006_),
    .B2(net161),
    .C1(_00025_),
    .X(_00040_));
 sky130_fd_sc_hd__a211o_1 _24377_ (.A1(_00009_),
    .A2(_00024_),
    .B1(_08296_),
    .C1(_08298_),
    .X(_00041_));
 sky130_fd_sc_hd__nand3_2 _24378_ (.A(_00036_),
    .B(_00030_),
    .C(_00034_),
    .Y(_00042_));
 sky130_fd_sc_hd__o22ai_4 _24379_ (.A1(_14098_),
    .A2(_00028_),
    .B1(_00032_),
    .B2(_00035_),
    .Y(_00043_));
 sky130_fd_sc_hd__nand3_2 _24380_ (.A(_00043_),
    .B(net159),
    .C(_00042_),
    .Y(_00045_));
 sky130_fd_sc_hd__a31oi_4 _24381_ (.A1(_00043_),
    .A2(net159),
    .A3(_00042_),
    .B1(_00040_),
    .Y(_00046_));
 sky130_fd_sc_hd__o211ai_4 _24382_ (.A1(_00026_),
    .A2(net159),
    .B1(_04238_),
    .C1(_00039_),
    .Y(_00047_));
 sky130_fd_sc_hd__and3_1 _24383_ (.A(_00045_),
    .B(_04227_),
    .C(_00041_),
    .X(_00048_));
 sky130_fd_sc_hd__nand3_2 _24384_ (.A(_00045_),
    .B(_04227_),
    .C(_00041_),
    .Y(_00049_));
 sky130_fd_sc_hd__o21a_1 _24385_ (.A1(_02137_),
    .A2(_14108_),
    .B1(_14115_),
    .X(_00050_));
 sky130_fd_sc_hd__o21ai_4 _24386_ (.A1(_14115_),
    .A2(_14112_),
    .B1(_14111_),
    .Y(_00051_));
 sky130_fd_sc_hd__a21oi_1 _24387_ (.A1(_14114_),
    .A2(_14113_),
    .B1(_14110_),
    .Y(_00052_));
 sky130_fd_sc_hd__or3_2 _24388_ (.A(net158),
    .B(_08712_),
    .C(_00046_),
    .X(_00053_));
 sky130_fd_sc_hd__a21oi_4 _24389_ (.A1(_00047_),
    .A2(_00049_),
    .B1(_00051_),
    .Y(_00054_));
 sky130_fd_sc_hd__o2bb2ai_1 _24390_ (.A1_N(_00047_),
    .A2_N(_00049_),
    .B1(_00050_),
    .B2(_14112_),
    .Y(_00056_));
 sky130_fd_sc_hd__nand3_1 _24391_ (.A(_00047_),
    .B(_00049_),
    .C(_00051_),
    .Y(_00057_));
 sky130_fd_sc_hd__a31o_2 _24392_ (.A1(_00047_),
    .A2(_00049_),
    .A3(_00051_),
    .B1(_08715_),
    .X(_00058_));
 sky130_fd_sc_hd__nand3_4 _24393_ (.A(_00056_),
    .B(_00057_),
    .C(_08714_),
    .Y(_00059_));
 sky130_fd_sc_hd__o22ai_4 _24394_ (.A1(_08714_),
    .A2(_00046_),
    .B1(_00054_),
    .B2(_00058_),
    .Y(_00060_));
 sky130_fd_sc_hd__a2bb2oi_4 _24395_ (.A1_N(_02049_),
    .A2_N(net343),
    .B1(_00053_),
    .B2(_00059_),
    .Y(_00061_));
 sky130_fd_sc_hd__o21ai_4 _24396_ (.A1(_02049_),
    .A2(net343),
    .B1(_00060_),
    .Y(_00062_));
 sky130_fd_sc_hd__o221a_2 _24397_ (.A1(_08714_),
    .A2(_00046_),
    .B1(_00054_),
    .B2(_00058_),
    .C1(_02137_),
    .X(_00063_));
 sky130_fd_sc_hd__o221ai_4 _24398_ (.A1(_08714_),
    .A2(_00046_),
    .B1(_00054_),
    .B2(_00058_),
    .C1(_02137_),
    .Y(_00064_));
 sky130_fd_sc_hd__and4_1 _24399_ (.A(_12793_),
    .B(_12795_),
    .C(_13271_),
    .D(_13274_),
    .X(_00065_));
 sky130_fd_sc_hd__nand3_1 _24400_ (.A(_14130_),
    .B(_00065_),
    .C(_13711_),
    .Y(_00067_));
 sky130_fd_sc_hd__o211ai_4 _24401_ (.A1(_14136_),
    .A2(_14128_),
    .B1(_14132_),
    .C1(_00067_),
    .Y(_00068_));
 sky130_fd_sc_hd__nor4b_1 _24402_ (.A(_12798_),
    .B(_13707_),
    .C(_13709_),
    .D_N(_00065_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand4_4 _24403_ (.A(_14130_),
    .B(_00065_),
    .C(_12797_),
    .D(_13711_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand3_1 _24404_ (.A(_00069_),
    .B(_14132_),
    .C(_14130_),
    .Y(_00071_));
 sky130_fd_sc_hd__o31a_1 _24405_ (.A1(_12798_),
    .A2(_14131_),
    .A3(_00067_),
    .B1(_00068_),
    .X(_00072_));
 sky130_fd_sc_hd__o21ai_4 _24406_ (.A1(_14131_),
    .A2(_00070_),
    .B1(_00068_),
    .Y(_00073_));
 sky130_fd_sc_hd__o21ai_4 _24407_ (.A1(_00061_),
    .A2(_00063_),
    .B1(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__o211ai_4 _24408_ (.A1(_00070_),
    .A2(_14131_),
    .B1(_00064_),
    .C1(_00068_),
    .Y(_00075_));
 sky130_fd_sc_hd__o2111ai_4 _24409_ (.A1(_14131_),
    .A2(_00070_),
    .B1(_00068_),
    .C1(_00064_),
    .D1(_00062_),
    .Y(_00076_));
 sky130_fd_sc_hd__o221ai_4 _24410_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_00061_),
    .B2(_00075_),
    .C1(_00074_),
    .Y(_00078_));
 sky130_fd_sc_hd__a21oi_2 _24411_ (.A1(_00053_),
    .A2(_00059_),
    .B1(_09125_),
    .Y(_00079_));
 sky130_fd_sc_hd__a211o_4 _24412_ (.A1(_00053_),
    .A2(_00059_),
    .B1(_09120_),
    .C1(_09121_),
    .X(_00080_));
 sky130_fd_sc_hd__a31oi_4 _24413_ (.A1(_09125_),
    .A2(_00074_),
    .A3(_00076_),
    .B1(_00079_),
    .Y(_00081_));
 sky130_fd_sc_hd__a21oi_4 _24414_ (.A1(_00078_),
    .A2(_00080_),
    .B1(net143),
    .Y(_00082_));
 sky130_fd_sc_hd__or3_1 _24415_ (.A(_09553_),
    .B(net155),
    .C(_00081_),
    .X(_00083_));
 sky130_fd_sc_hd__a311oi_4 _24416_ (.A1(_09125_),
    .A2(_00074_),
    .A3(_00076_),
    .B1(_00079_),
    .C1(_00251_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand3_2 _24417_ (.A(_00078_),
    .B(_00080_),
    .C(_00240_),
    .Y(_00085_));
 sky130_fd_sc_hd__a22oi_4 _24418_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_00078_),
    .B2(_00080_),
    .Y(_00086_));
 sky130_fd_sc_hd__a22o_2 _24419_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_00078_),
    .B2(_00080_),
    .X(_00087_));
 sky130_fd_sc_hd__o22a_1 _24420_ (.A1(_14149_),
    .A2(_14126_),
    .B1(_14148_),
    .B2(_14152_),
    .X(_00089_));
 sky130_fd_sc_hd__o22ai_4 _24421_ (.A1(_14149_),
    .A2(_14126_),
    .B1(_14148_),
    .B2(_14152_),
    .Y(_00090_));
 sky130_fd_sc_hd__o21ai_4 _24422_ (.A1(_00084_),
    .A2(_00086_),
    .B1(_00090_),
    .Y(_00091_));
 sky130_fd_sc_hd__nand3_4 _24423_ (.A(_00085_),
    .B(_00087_),
    .C(_00089_),
    .Y(_00092_));
 sky130_fd_sc_hd__o311ai_4 _24424_ (.A1(_00084_),
    .A2(_00090_),
    .A3(_00086_),
    .B1(net143),
    .C1(_00091_),
    .Y(_00093_));
 sky130_fd_sc_hd__a31oi_4 _24425_ (.A1(net143),
    .A2(_00091_),
    .A3(_00092_),
    .B1(_00082_),
    .Y(_00094_));
 sky130_fd_sc_hd__a31o_1 _24426_ (.A1(net143),
    .A2(_00091_),
    .A3(_00092_),
    .B1(_00082_),
    .X(_00095_));
 sky130_fd_sc_hd__a311o_1 _24427_ (.A1(net143),
    .A2(_00091_),
    .A3(_00092_),
    .B1(_09579_),
    .C1(_00082_),
    .X(_00096_));
 sky130_fd_sc_hd__and3_1 _24428_ (.A(_13741_),
    .B(_13751_),
    .C(_14161_),
    .X(_00097_));
 sky130_fd_sc_hd__o21ai_2 _24429_ (.A1(_14166_),
    .A2(_14163_),
    .B1(_14161_),
    .Y(_00098_));
 sky130_fd_sc_hd__a311oi_4 _24430_ (.A1(net143),
    .A2(_00091_),
    .A3(_00092_),
    .B1(_00082_),
    .C1(_12899_),
    .Y(_00099_));
 sky130_fd_sc_hd__o221ai_4 _24431_ (.A1(_12867_),
    .A2(_12877_),
    .B1(net143),
    .B2(_00081_),
    .C1(_00093_),
    .Y(_00100_));
 sky130_fd_sc_hd__a21oi_2 _24432_ (.A1(_00083_),
    .A2(_00093_),
    .B1(_12888_),
    .Y(_00101_));
 sky130_fd_sc_hd__a2bb2o_1 _24433_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_00083_),
    .B2(_00093_),
    .X(_00102_));
 sky130_fd_sc_hd__o211ai_1 _24434_ (.A1(_14163_),
    .A2(_00097_),
    .B1(_00100_),
    .C1(_00102_),
    .Y(_00103_));
 sky130_fd_sc_hd__o21ai_1 _24435_ (.A1(_00099_),
    .A2(_00101_),
    .B1(_00098_),
    .Y(_00104_));
 sky130_fd_sc_hd__o211ai_2 _24436_ (.A1(_09571_),
    .A2(_09573_),
    .B1(_00103_),
    .C1(_00104_),
    .Y(_00105_));
 sky130_fd_sc_hd__o21ai_1 _24437_ (.A1(_12888_),
    .A2(_00094_),
    .B1(_00098_),
    .Y(_00106_));
 sky130_fd_sc_hd__o22ai_1 _24438_ (.A1(_14163_),
    .A2(_00097_),
    .B1(_00099_),
    .B2(_00101_),
    .Y(_00107_));
 sky130_fd_sc_hd__o211ai_2 _24439_ (.A1(_00099_),
    .A2(_00106_),
    .B1(_00107_),
    .C1(_09579_),
    .Y(_00108_));
 sky130_fd_sc_hd__o21ai_1 _24440_ (.A1(_09579_),
    .A2(_00094_),
    .B1(_00108_),
    .Y(_00110_));
 sky130_fd_sc_hd__inv_2 _24441_ (.A(_00110_),
    .Y(_00111_));
 sky130_fd_sc_hd__o211ai_4 _24442_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_00096_),
    .C1(_00105_),
    .Y(_00112_));
 sky130_fd_sc_hd__o211a_1 _24443_ (.A1(_09579_),
    .A2(_00094_),
    .B1(_11298_),
    .C1(_00108_),
    .X(_00113_));
 sky130_fd_sc_hd__o211ai_2 _24444_ (.A1(_09579_),
    .A2(_00094_),
    .B1(_11298_),
    .C1(_00108_),
    .Y(_00114_));
 sky130_fd_sc_hd__o32a_1 _24445_ (.A1(_10025_),
    .A2(_14167_),
    .A3(_14170_),
    .B1(_14179_),
    .B2(_14174_),
    .X(_00115_));
 sky130_fd_sc_hd__a21oi_2 _24446_ (.A1(_00112_),
    .A2(_00114_),
    .B1(_00115_),
    .Y(_00116_));
 sky130_fd_sc_hd__a31o_1 _24447_ (.A1(_00112_),
    .A2(_00115_),
    .A3(_00114_),
    .B1(_10479_),
    .X(_00117_));
 sky130_fd_sc_hd__o22ai_1 _24448_ (.A1(_10480_),
    .A2(_00111_),
    .B1(_00116_),
    .B2(_00117_),
    .Y(_00118_));
 sky130_fd_sc_hd__o221a_1 _24449_ (.A1(_10480_),
    .A2(_00111_),
    .B1(_00116_),
    .B2(_00117_),
    .C1(_10953_),
    .X(_00119_));
 sky130_fd_sc_hd__o21ai_2 _24450_ (.A1(_09927_),
    .A2(_09949_),
    .B1(_00118_),
    .Y(_00121_));
 sky130_fd_sc_hd__o221a_1 _24451_ (.A1(net131),
    .A2(_00111_),
    .B1(_00116_),
    .B2(_00117_),
    .C1(_10015_),
    .X(_00122_));
 sky130_fd_sc_hd__o221ai_4 _24452_ (.A1(_10480_),
    .A2(_00111_),
    .B1(_00116_),
    .B2(_00117_),
    .C1(_10015_),
    .Y(_00123_));
 sky130_fd_sc_hd__a21boi_2 _24453_ (.A1(_14188_),
    .A2(_14189_),
    .B1_N(_14190_),
    .Y(_00124_));
 sky130_fd_sc_hd__nand3_1 _24454_ (.A(_00121_),
    .B(_00123_),
    .C(_00124_),
    .Y(_00125_));
 sky130_fd_sc_hd__a21o_1 _24455_ (.A1(_00121_),
    .A2(_00123_),
    .B1(_00124_),
    .X(_00126_));
 sky130_fd_sc_hd__a31oi_2 _24456_ (.A1(_10954_),
    .A2(_00125_),
    .A3(_00126_),
    .B1(_00119_),
    .Y(_00127_));
 sky130_fd_sc_hd__a21oi_1 _24457_ (.A1(_07899_),
    .A2(_14193_),
    .B1(_14200_),
    .Y(_00128_));
 sky130_fd_sc_hd__a21oi_1 _24458_ (.A1(_08874_),
    .A2(_08896_),
    .B1(_00127_),
    .Y(_00129_));
 sky130_fd_sc_hd__or3_1 _24459_ (.A(_08819_),
    .B(_08841_),
    .C(_00127_),
    .X(_00130_));
 sky130_fd_sc_hd__a311o_1 _24460_ (.A1(_10954_),
    .A2(_00125_),
    .A3(_00126_),
    .B1(_00119_),
    .C1(_08907_),
    .X(_00132_));
 sky130_fd_sc_hd__a21oi_1 _24461_ (.A1(_00130_),
    .A2(_00132_),
    .B1(_00128_),
    .Y(_00133_));
 sky130_fd_sc_hd__a31o_1 _24462_ (.A1(_00130_),
    .A2(_00132_),
    .A3(_00128_),
    .B1(_11464_),
    .X(_00134_));
 sky130_fd_sc_hd__o22ai_2 _24463_ (.A1(_11465_),
    .A2(_00127_),
    .B1(_00133_),
    .B2(_00134_),
    .Y(_00135_));
 sky130_fd_sc_hd__o21bai_1 _24464_ (.A1(_14204_),
    .A2(_14205_),
    .B1_N(_14203_),
    .Y(_00136_));
 sky130_fd_sc_hd__o21ai_1 _24465_ (.A1(net368),
    .A2(_07866_),
    .B1(_00135_),
    .Y(_00137_));
 sky130_fd_sc_hd__o221a_1 _24466_ (.A1(_11465_),
    .A2(_00127_),
    .B1(_00133_),
    .B2(_00134_),
    .C1(_07899_),
    .X(_00138_));
 sky130_fd_sc_hd__or3_1 _24467_ (.A(net368),
    .B(_07866_),
    .C(_00135_),
    .X(_00139_));
 sky130_fd_sc_hd__a21oi_1 _24468_ (.A1(_00137_),
    .A2(_00139_),
    .B1(_00136_),
    .Y(_00140_));
 sky130_fd_sc_hd__o21ai_1 _24469_ (.A1(_11944_),
    .A2(_00140_),
    .B1(_00135_),
    .Y(_00141_));
 sky130_fd_sc_hd__or3_1 _24470_ (.A(_05051_),
    .B(_14209_),
    .C(_00141_),
    .X(_00143_));
 sky130_fd_sc_hd__o21ai_1 _24471_ (.A1(_05051_),
    .A2(_14209_),
    .B1(_00141_),
    .Y(_00144_));
 sky130_fd_sc_hd__nand2_1 _24472_ (.A(_00143_),
    .B(_00144_),
    .Y(net95));
 sky130_fd_sc_hd__o211ai_1 _24473_ (.A1(_11944_),
    .A2(_00140_),
    .B1(_00135_),
    .C1(_14209_),
    .Y(_00145_));
 sky130_fd_sc_hd__o211ai_2 _24474_ (.A1(_14211_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_14220_),
    .Y(_00146_));
 sky130_fd_sc_hd__and3_1 _24475_ (.A(_00146_),
    .B(net335),
    .C(_11079_),
    .X(_00147_));
 sky130_fd_sc_hd__a311o_2 _24476_ (.A1(_11471_),
    .A2(_14213_),
    .A3(_14220_),
    .B1(net332),
    .C1(_09840_),
    .X(_00148_));
 sky130_fd_sc_hd__o211ai_2 _24477_ (.A1(net351),
    .A2(_09807_),
    .B1(_10971_),
    .C1(_00146_),
    .Y(_00149_));
 sky130_fd_sc_hd__o2bb2ai_1 _24478_ (.A1_N(net335),
    .A2_N(_00146_),
    .B1(_10967_),
    .B2(_10965_),
    .Y(_00150_));
 sky130_fd_sc_hd__and2_1 _24479_ (.A(_00149_),
    .B(_00150_),
    .X(_00151_));
 sky130_fd_sc_hd__nand2_1 _24480_ (.A(_00149_),
    .B(_00150_),
    .Y(_00153_));
 sky130_fd_sc_hd__o21ai_2 _24481_ (.A1(_14229_),
    .A2(_14232_),
    .B1(_14228_),
    .Y(_00154_));
 sky130_fd_sc_hd__nand2_2 _24482_ (.A(_00154_),
    .B(_00151_),
    .Y(_00155_));
 sky130_fd_sc_hd__o211ai_1 _24483_ (.A1(_14229_),
    .A2(_14232_),
    .B1(_00153_),
    .C1(_14228_),
    .Y(_00156_));
 sky130_fd_sc_hd__o221ai_4 _24484_ (.A1(_11046_),
    .A2(_11057_),
    .B1(_00151_),
    .B2(_00154_),
    .C1(_00155_),
    .Y(_00157_));
 sky130_fd_sc_hd__a21oi_4 _24485_ (.A1(_00148_),
    .A2(_00157_),
    .B1(net311),
    .Y(_00158_));
 sky130_fd_sc_hd__a21oi_1 _24486_ (.A1(_00148_),
    .A2(_00157_),
    .B1(net150),
    .Y(_00159_));
 sky130_fd_sc_hd__a2bb2o_2 _24487_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_00148_),
    .B2(_00157_),
    .X(_00160_));
 sky130_fd_sc_hd__a31o_1 _24488_ (.A1(_00155_),
    .A2(_00156_),
    .A3(net332),
    .B1(_10492_),
    .X(_00161_));
 sky130_fd_sc_hd__and3_1 _24489_ (.A(_00157_),
    .B(net150),
    .C(_00148_),
    .X(_00162_));
 sky130_fd_sc_hd__o21ai_2 _24490_ (.A1(_00147_),
    .A2(_00161_),
    .B1(_00160_),
    .Y(_00164_));
 sky130_fd_sc_hd__a31oi_4 _24491_ (.A1(_14242_),
    .A2(_14245_),
    .A3(_14247_),
    .B1(_14240_),
    .Y(_00165_));
 sky130_fd_sc_hd__a31o_1 _24492_ (.A1(_14242_),
    .A2(_14245_),
    .A3(_14247_),
    .B1(_14240_),
    .X(_00166_));
 sky130_fd_sc_hd__o21ai_2 _24493_ (.A1(_00159_),
    .A2(_00162_),
    .B1(_00165_),
    .Y(_00167_));
 sky130_fd_sc_hd__o211ai_1 _24494_ (.A1(_00161_),
    .A2(_00147_),
    .B1(_00160_),
    .C1(_00166_),
    .Y(_00168_));
 sky130_fd_sc_hd__o221a_2 _24495_ (.A1(net329),
    .A2(net327),
    .B1(_00165_),
    .B2(_00164_),
    .C1(_00167_),
    .X(_00169_));
 sky130_fd_sc_hd__o221ai_4 _24496_ (.A1(net329),
    .A2(net327),
    .B1(_00165_),
    .B2(_00164_),
    .C1(_00167_),
    .Y(_00170_));
 sky130_fd_sc_hd__nor2_2 _24497_ (.A(_00158_),
    .B(_00169_),
    .Y(_00171_));
 sky130_fd_sc_hd__o22a_1 _24498_ (.A1(_14458_),
    .A2(_00000_),
    .B1(_00158_),
    .B2(_00169_),
    .X(_00172_));
 sky130_fd_sc_hd__or3_1 _24499_ (.A(_00011_),
    .B(net323),
    .C(_00171_),
    .X(_00173_));
 sky130_fd_sc_hd__o22a_1 _24500_ (.A1(net170),
    .A2(net169),
    .B1(_00158_),
    .B2(_00169_),
    .X(_00175_));
 sky130_fd_sc_hd__o22ai_4 _24501_ (.A1(net170),
    .A2(net169),
    .B1(_00158_),
    .B2(_00169_),
    .Y(_00176_));
 sky130_fd_sc_hd__nand3b_4 _24502_ (.A_N(_00158_),
    .B(_00170_),
    .C(net153),
    .Y(_00177_));
 sky130_fd_sc_hd__nand2_1 _24503_ (.A(_00176_),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__and3_1 _24504_ (.A(_12985_),
    .B(_13413_),
    .C(_13414_),
    .X(_00179_));
 sky130_fd_sc_hd__nand3_1 _24505_ (.A(_14262_),
    .B(_00179_),
    .C(_13859_),
    .Y(_00180_));
 sky130_fd_sc_hd__o211ai_4 _24506_ (.A1(_14259_),
    .A2(_14261_),
    .B1(_14264_),
    .C1(_00180_),
    .Y(_00181_));
 sky130_fd_sc_hd__nor4b_1 _24507_ (.A(_12994_),
    .B(_13855_),
    .C(_13857_),
    .D_N(_00179_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand3_4 _24508_ (.A(_00182_),
    .B(_14264_),
    .C(_14262_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand2_1 _24509_ (.A(_00181_),
    .B(_00183_),
    .Y(_00184_));
 sky130_fd_sc_hd__a22oi_1 _24510_ (.A1(_00176_),
    .A2(_00177_),
    .B1(_00181_),
    .B2(_00183_),
    .Y(_00186_));
 sky130_fd_sc_hd__a22o_1 _24511_ (.A1(_00176_),
    .A2(_00177_),
    .B1(_00181_),
    .B2(_00183_),
    .X(_00187_));
 sky130_fd_sc_hd__nand4_4 _24512_ (.A(_00176_),
    .B(_00177_),
    .C(_00181_),
    .D(_00183_),
    .Y(_00188_));
 sky130_fd_sc_hd__o22ai_1 _24513_ (.A1(_00011_),
    .A2(net321),
    .B1(_00178_),
    .B2(_00184_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand3_4 _24514_ (.A(_00187_),
    .B(_00188_),
    .C(net308),
    .Y(_00190_));
 sky130_fd_sc_hd__o22ai_2 _24515_ (.A1(net308),
    .A2(_00171_),
    .B1(_00186_),
    .B2(_00189_),
    .Y(_00191_));
 sky130_fd_sc_hd__a21oi_2 _24516_ (.A1(_00173_),
    .A2(_00190_),
    .B1(net278),
    .Y(_00192_));
 sky130_fd_sc_hd__a211o_1 _24517_ (.A1(_00173_),
    .A2(_00190_),
    .B1(net304),
    .C1(_01951_),
    .X(_00193_));
 sky130_fd_sc_hd__a311oi_4 _24518_ (.A1(_00187_),
    .A2(_00188_),
    .A3(net308),
    .B1(_09595_),
    .C1(_00172_),
    .Y(_00194_));
 sky130_fd_sc_hd__o211ai_4 _24519_ (.A1(net307),
    .A2(_00171_),
    .B1(net172),
    .C1(_00190_),
    .Y(_00195_));
 sky130_fd_sc_hd__a22oi_1 _24520_ (.A1(_09589_),
    .A2(_09591_),
    .B1(_00173_),
    .B2(_00190_),
    .Y(_00197_));
 sky130_fd_sc_hd__o21ai_4 _24521_ (.A1(_09588_),
    .A2(_09590_),
    .B1(_00191_),
    .Y(_00198_));
 sky130_fd_sc_hd__a31o_1 _24522_ (.A1(_13871_),
    .A2(_14272_),
    .A3(_14276_),
    .B1(_14273_),
    .X(_00199_));
 sky130_fd_sc_hd__a31oi_4 _24523_ (.A1(_13871_),
    .A2(_14272_),
    .A3(_14276_),
    .B1(_14273_),
    .Y(_00200_));
 sky130_fd_sc_hd__o21ai_2 _24524_ (.A1(_00194_),
    .A2(_00197_),
    .B1(_00200_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand3_2 _24525_ (.A(_00195_),
    .B(_00198_),
    .C(_00199_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand3_1 _24526_ (.A(_00201_),
    .B(_00202_),
    .C(net278),
    .Y(_00203_));
 sky130_fd_sc_hd__a31oi_1 _24527_ (.A1(_00201_),
    .A2(_00202_),
    .A3(net278),
    .B1(_00192_),
    .Y(_00204_));
 sky130_fd_sc_hd__a31o_1 _24528_ (.A1(_00201_),
    .A2(_00202_),
    .A3(net278),
    .B1(_00192_),
    .X(_00205_));
 sky130_fd_sc_hd__a21boi_1 _24529_ (.A1(_14291_),
    .A2(_14287_),
    .B1_N(_14286_),
    .Y(_00206_));
 sky130_fd_sc_hd__o22ai_4 _24530_ (.A1(net177),
    .A2(_14285_),
    .B1(_14288_),
    .B2(_14292_),
    .Y(_00208_));
 sky130_fd_sc_hd__a311oi_2 _24531_ (.A1(_00201_),
    .A2(_00202_),
    .A3(net278),
    .B1(net173),
    .C1(_00192_),
    .Y(_00209_));
 sky130_fd_sc_hd__a311o_1 _24532_ (.A1(_00201_),
    .A2(_00202_),
    .A3(net278),
    .B1(net173),
    .C1(_00192_),
    .X(_00210_));
 sky130_fd_sc_hd__a2bb2oi_2 _24533_ (.A1_N(_09134_),
    .A2_N(_09135_),
    .B1(_00193_),
    .B2(_00203_),
    .Y(_00211_));
 sky130_fd_sc_hd__a2bb2o_1 _24534_ (.A1_N(_09134_),
    .A2_N(_09135_),
    .B1(_00193_),
    .B2(_00203_),
    .X(_00212_));
 sky130_fd_sc_hd__nor2_1 _24535_ (.A(_00209_),
    .B(_00211_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand3_2 _24536_ (.A(_00208_),
    .B(_00210_),
    .C(_00212_),
    .Y(_00214_));
 sky130_fd_sc_hd__o21ai_2 _24537_ (.A1(_00209_),
    .A2(_00211_),
    .B1(_00206_),
    .Y(_00215_));
 sky130_fd_sc_hd__a21oi_2 _24538_ (.A1(_00193_),
    .A2(_00203_),
    .B1(_04029_),
    .Y(_00216_));
 sky130_fd_sc_hd__or3_1 _24539_ (.A(net302),
    .B(_04019_),
    .C(_00204_),
    .X(_00217_));
 sky130_fd_sc_hd__nand3_2 _24540_ (.A(_00214_),
    .B(_00215_),
    .C(_04029_),
    .Y(_00219_));
 sky130_fd_sc_hd__a31oi_4 _24541_ (.A1(_00214_),
    .A2(_00215_),
    .A3(_04029_),
    .B1(_00216_),
    .Y(_00220_));
 sky130_fd_sc_hd__a2bb2oi_1 _24542_ (.A1_N(_08724_),
    .A2_N(net196),
    .B1(_00217_),
    .B2(_00219_),
    .Y(_00221_));
 sky130_fd_sc_hd__a22o_1 _24543_ (.A1(_08725_),
    .A2(_08727_),
    .B1(_00217_),
    .B2(_00219_),
    .X(_00222_));
 sky130_fd_sc_hd__o211a_1 _24544_ (.A1(_04029_),
    .A2(_00204_),
    .B1(net177),
    .C1(_00219_),
    .X(_00223_));
 sky130_fd_sc_hd__a311o_1 _24545_ (.A1(_00214_),
    .A2(_00215_),
    .A3(_04029_),
    .B1(_00216_),
    .C1(net175),
    .X(_00224_));
 sky130_fd_sc_hd__nand2_1 _24546_ (.A(_14310_),
    .B(_14316_),
    .Y(_00225_));
 sky130_fd_sc_hd__o211ai_1 _24547_ (.A1(_14300_),
    .A2(net198),
    .B1(_14310_),
    .C1(_14309_),
    .Y(_00226_));
 sky130_fd_sc_hd__o22ai_1 _24548_ (.A1(net199),
    .A2(_14301_),
    .B1(_00225_),
    .B2(_14308_),
    .Y(_00227_));
 sky130_fd_sc_hd__a31oi_2 _24549_ (.A1(_14309_),
    .A2(_14310_),
    .A3(_14316_),
    .B1(_14312_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand3_2 _24550_ (.A(_00227_),
    .B(_00224_),
    .C(_00222_),
    .Y(_00230_));
 sky130_fd_sc_hd__o21ai_2 _24551_ (.A1(_00221_),
    .A2(_00223_),
    .B1(_00228_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand3_1 _24552_ (.A(_00230_),
    .B(_00231_),
    .C(net271),
    .Y(_00232_));
 sky130_fd_sc_hd__a21oi_2 _24553_ (.A1(_00217_),
    .A2(_00219_),
    .B1(net271),
    .Y(_00233_));
 sky130_fd_sc_hd__or3_1 _24554_ (.A(net296),
    .B(_05232_),
    .C(_00220_),
    .X(_00234_));
 sky130_fd_sc_hd__o31a_2 _24555_ (.A1(net296),
    .A2(_05232_),
    .A3(_00220_),
    .B1(_00232_),
    .X(_00235_));
 sky130_fd_sc_hd__a31o_1 _24556_ (.A1(_00230_),
    .A2(_00231_),
    .A3(net271),
    .B1(_00233_),
    .X(_00236_));
 sky130_fd_sc_hd__a311o_1 _24557_ (.A1(_00230_),
    .A2(_00231_),
    .A3(net271),
    .B1(_00233_),
    .C1(net244),
    .X(_00237_));
 sky130_fd_sc_hd__a22oi_2 _24558_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_00232_),
    .B2(_00234_),
    .Y(_00238_));
 sky130_fd_sc_hd__a22o_1 _24559_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_00232_),
    .B2(_00234_),
    .X(_00239_));
 sky130_fd_sc_hd__a31oi_1 _24560_ (.A1(_00230_),
    .A2(_00231_),
    .A3(net271),
    .B1(net198),
    .Y(_00241_));
 sky130_fd_sc_hd__a31o_1 _24561_ (.A1(_00230_),
    .A2(_00231_),
    .A3(net271),
    .B1(net198),
    .X(_00242_));
 sky130_fd_sc_hd__and3_1 _24562_ (.A(_00232_),
    .B(_00234_),
    .C(net199),
    .X(_00243_));
 sky130_fd_sc_hd__a311o_1 _24563_ (.A1(_00230_),
    .A2(_00231_),
    .A3(net271),
    .B1(_00233_),
    .C1(net198),
    .X(_00244_));
 sky130_fd_sc_hd__a21oi_1 _24564_ (.A1(_00234_),
    .A2(_00241_),
    .B1(_00238_),
    .Y(_00245_));
 sky130_fd_sc_hd__and3_1 _24565_ (.A(_13060_),
    .B(_13486_),
    .C(_13488_),
    .X(_00246_));
 sky130_fd_sc_hd__nor4_1 _24566_ (.A(_13061_),
    .B(_13489_),
    .C(_13932_),
    .D(_13934_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand3_1 _24567_ (.A(_14329_),
    .B(_00246_),
    .C(_13936_),
    .Y(_00248_));
 sky130_fd_sc_hd__o211ai_4 _24568_ (.A1(_14333_),
    .A2(_14328_),
    .B1(_14331_),
    .C1(_00248_),
    .Y(_00249_));
 sky130_fd_sc_hd__o2111a_1 _24569_ (.A1(_13068_),
    .A2(_13073_),
    .B1(_13933_),
    .C1(_00246_),
    .D1(_13935_),
    .X(_00250_));
 sky130_fd_sc_hd__o211ai_2 _24570_ (.A1(_07935_),
    .A2(_14323_),
    .B1(_13076_),
    .C1(_00247_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand3_4 _24571_ (.A(_14329_),
    .B(_14331_),
    .C(_00250_),
    .Y(_00253_));
 sky130_fd_sc_hd__o21ai_4 _24572_ (.A1(_14328_),
    .A2(_00252_),
    .B1(_00249_),
    .Y(_00254_));
 sky130_fd_sc_hd__inv_2 _24573_ (.A(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _24574_ (.A(_00254_),
    .B(_00245_),
    .Y(_00256_));
 sky130_fd_sc_hd__o211ai_1 _24575_ (.A1(_00238_),
    .A2(_00243_),
    .B1(_00249_),
    .C1(_00253_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand4_2 _24576_ (.A(_00239_),
    .B(_00244_),
    .C(_00249_),
    .D(_00253_),
    .Y(_00258_));
 sky130_fd_sc_hd__o21ai_2 _24577_ (.A1(_00238_),
    .A2(_00243_),
    .B1(_00254_),
    .Y(_00259_));
 sky130_fd_sc_hd__nand3_2 _24578_ (.A(_00256_),
    .B(_00257_),
    .C(net244),
    .Y(_00260_));
 sky130_fd_sc_hd__and3_1 _24579_ (.A(_05482_),
    .B(_05484_),
    .C(_00236_),
    .X(_00261_));
 sky130_fd_sc_hd__inv_2 _24580_ (.A(_00261_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand3_2 _24581_ (.A(_00259_),
    .B(net244),
    .C(_00258_),
    .Y(_00264_));
 sky130_fd_sc_hd__and3_2 _24582_ (.A(_05754_),
    .B(_00237_),
    .C(_00260_),
    .X(_00265_));
 sky130_fd_sc_hd__a211o_2 _24583_ (.A1(_00263_),
    .A2(_00264_),
    .B1(net265),
    .C1(net264),
    .X(_00266_));
 sky130_fd_sc_hd__a311oi_4 _24584_ (.A1(_00259_),
    .A2(net244),
    .A3(_00258_),
    .B1(_00261_),
    .C1(_07936_),
    .Y(_00267_));
 sky130_fd_sc_hd__nand3_4 _24585_ (.A(_00264_),
    .B(_07935_),
    .C(_00263_),
    .Y(_00268_));
 sky130_fd_sc_hd__o211ai_4 _24586_ (.A1(_00236_),
    .A2(net244),
    .B1(_07936_),
    .C1(_00260_),
    .Y(_00269_));
 sky130_fd_sc_hd__a21oi_1 _24587_ (.A1(_13948_),
    .A2(_14340_),
    .B1(_14345_),
    .Y(_00270_));
 sky130_fd_sc_hd__a31o_1 _24588_ (.A1(_13948_),
    .A2(_14340_),
    .A3(_14344_),
    .B1(_14345_),
    .X(_00271_));
 sky130_fd_sc_hd__a31oi_4 _24589_ (.A1(_13948_),
    .A2(_14340_),
    .A3(_14344_),
    .B1(_14345_),
    .Y(_00272_));
 sky130_fd_sc_hd__o2bb2ai_4 _24590_ (.A1_N(_00268_),
    .A2_N(_00269_),
    .B1(_00270_),
    .B2(_14343_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand3_4 _24591_ (.A(_00271_),
    .B(_00269_),
    .C(_00268_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand3_2 _24592_ (.A(_00274_),
    .B(_00275_),
    .C(net243),
    .Y(_00276_));
 sky130_fd_sc_hd__a31oi_4 _24593_ (.A1(_00274_),
    .A2(_00275_),
    .A3(net243),
    .B1(_00265_),
    .Y(_00277_));
 sky130_fd_sc_hd__a311o_1 _24594_ (.A1(_00274_),
    .A2(_00275_),
    .A3(net243),
    .B1(net240),
    .C1(_00265_),
    .X(_00278_));
 sky130_fd_sc_hd__o211ai_4 _24595_ (.A1(net227),
    .A2(_13960_),
    .B1(_14360_),
    .C1(_14365_),
    .Y(_00279_));
 sky130_fd_sc_hd__a31o_1 _24596_ (.A1(_13973_),
    .A2(_14360_),
    .A3(_14365_),
    .B1(_14361_),
    .X(_00280_));
 sky130_fd_sc_hd__a31oi_2 _24597_ (.A1(_00274_),
    .A2(_00275_),
    .A3(net243),
    .B1(net202),
    .Y(_00281_));
 sky130_fd_sc_hd__a311oi_4 _24598_ (.A1(_00274_),
    .A2(_00275_),
    .A3(net243),
    .B1(net202),
    .C1(_00265_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand3_2 _24599_ (.A(_00276_),
    .B(_07564_),
    .C(_00266_),
    .Y(_00283_));
 sky130_fd_sc_hd__a2bb2oi_4 _24600_ (.A1_N(net221),
    .A2_N(net220),
    .B1(_00266_),
    .B2(_00276_),
    .Y(_00285_));
 sky130_fd_sc_hd__a22o_1 _24601_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_00266_),
    .B2(_00276_),
    .X(_00286_));
 sky130_fd_sc_hd__o2111ai_1 _24602_ (.A1(_14361_),
    .A2(_14366_),
    .B1(_00283_),
    .C1(_00286_),
    .D1(_14360_),
    .Y(_00287_));
 sky130_fd_sc_hd__o221ai_1 _24603_ (.A1(net223),
    .A2(_14356_),
    .B1(_00282_),
    .B2(_00285_),
    .C1(_00279_),
    .Y(_00288_));
 sky130_fd_sc_hd__o211ai_1 _24604_ (.A1(net260),
    .A2(net258),
    .B1(_00287_),
    .C1(_00288_),
    .Y(_00289_));
 sky130_fd_sc_hd__o221ai_4 _24605_ (.A1(_14356_),
    .A2(net223),
    .B1(_07564_),
    .B2(_00277_),
    .C1(_00279_),
    .Y(_00290_));
 sky130_fd_sc_hd__o21ai_1 _24606_ (.A1(_00282_),
    .A2(_00285_),
    .B1(_00280_),
    .Y(_00291_));
 sky130_fd_sc_hd__o221ai_4 _24607_ (.A1(net260),
    .A2(net258),
    .B1(_00282_),
    .B2(_00290_),
    .C1(_00291_),
    .Y(_00292_));
 sky130_fd_sc_hd__o21ai_4 _24608_ (.A1(net240),
    .A2(_00277_),
    .B1(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__o31a_2 _24609_ (.A1(net260),
    .A2(net258),
    .A3(_00277_),
    .B1(_00292_),
    .X(_00294_));
 sky130_fd_sc_hd__o211ai_2 _24610_ (.A1(_07242_),
    .A2(net248),
    .B1(_00278_),
    .C1(_00289_),
    .Y(_00296_));
 sky130_fd_sc_hd__o211ai_4 _24611_ (.A1(net240),
    .A2(_00277_),
    .B1(_07246_),
    .C1(_00292_),
    .Y(_00297_));
 sky130_fd_sc_hd__nand2_1 _24612_ (.A(_00296_),
    .B(_00297_),
    .Y(_00298_));
 sky130_fd_sc_hd__a31o_1 _24613_ (.A1(_14379_),
    .A2(_14384_),
    .A3(_14386_),
    .B1(_14376_),
    .X(_00299_));
 sky130_fd_sc_hd__a31oi_1 _24614_ (.A1(_14379_),
    .A2(_14384_),
    .A3(_14386_),
    .B1(_14376_),
    .Y(_00300_));
 sky130_fd_sc_hd__and4_1 _24615_ (.A(_14377_),
    .B(_14394_),
    .C(_00296_),
    .D(_00297_),
    .X(_00301_));
 sky130_fd_sc_hd__o2bb2ai_2 _24616_ (.A1_N(_00298_),
    .A2_N(_00299_),
    .B1(net239),
    .B2(_06292_),
    .Y(_00302_));
 sky130_fd_sc_hd__and3_1 _24617_ (.A(_06294_),
    .B(_00278_),
    .C(_00289_),
    .X(_00303_));
 sky130_fd_sc_hd__o311a_1 _24618_ (.A1(_06918_),
    .A2(_06920_),
    .A3(_14375_),
    .B1(_14394_),
    .C1(_00298_),
    .X(_00304_));
 sky130_fd_sc_hd__o21ai_2 _24619_ (.A1(_00298_),
    .A2(_00300_),
    .B1(net214),
    .Y(_00305_));
 sky130_fd_sc_hd__o22a_2 _24620_ (.A1(net214),
    .A2(_00293_),
    .B1(_00301_),
    .B2(_00302_),
    .X(_00307_));
 sky130_fd_sc_hd__o22a_2 _24621_ (.A1(net214),
    .A2(_00294_),
    .B1(_00304_),
    .B2(_00305_),
    .X(_00308_));
 sky130_fd_sc_hd__o221ai_4 _24622_ (.A1(net214),
    .A2(_00293_),
    .B1(_00301_),
    .B2(_00302_),
    .C1(_06924_),
    .Y(_00309_));
 sky130_fd_sc_hd__o21ai_1 _24623_ (.A1(_00304_),
    .A2(_00305_),
    .B1(net227),
    .Y(_00310_));
 sky130_fd_sc_hd__o221ai_4 _24624_ (.A1(net214),
    .A2(_00294_),
    .B1(_00304_),
    .B2(_00305_),
    .C1(net227),
    .Y(_00311_));
 sky130_fd_sc_hd__and4_1 _24625_ (.A(_13143_),
    .B(_13144_),
    .C(_13568_),
    .D(_13571_),
    .X(_00312_));
 sky130_fd_sc_hd__and3_1 _24626_ (.A(_14010_),
    .B(_14012_),
    .C(_00312_),
    .X(_00313_));
 sky130_fd_sc_hd__nand3_1 _24627_ (.A(_14400_),
    .B(_00312_),
    .C(_14013_),
    .Y(_00314_));
 sky130_fd_sc_hd__o211ai_4 _24628_ (.A1(_14405_),
    .A2(_14399_),
    .B1(_14401_),
    .C1(_00314_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand4_4 _24629_ (.A(_00313_),
    .B(_14401_),
    .C(_14400_),
    .D(_13151_),
    .Y(_00316_));
 sky130_fd_sc_hd__and2_1 _24630_ (.A(_00315_),
    .B(_00316_),
    .X(_00318_));
 sky130_fd_sc_hd__a22o_2 _24631_ (.A1(_00309_),
    .A2(_00311_),
    .B1(_00315_),
    .B2(_00316_),
    .X(_00319_));
 sky130_fd_sc_hd__nand3_2 _24632_ (.A(_00311_),
    .B(_00315_),
    .C(_00316_),
    .Y(_00320_));
 sky130_fd_sc_hd__o2111ai_4 _24633_ (.A1(_06924_),
    .A2(_00307_),
    .B1(_00309_),
    .C1(_00315_),
    .D1(_00316_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand3_2 _24634_ (.A(_00319_),
    .B(_00321_),
    .C(net210),
    .Y(_00322_));
 sky130_fd_sc_hd__o221a_2 _24635_ (.A1(net214),
    .A2(_00293_),
    .B1(_00301_),
    .B2(_00302_),
    .C1(_06613_),
    .X(_00323_));
 sky130_fd_sc_hd__or3_2 _24636_ (.A(net238),
    .B(_06610_),
    .C(_00308_),
    .X(_00324_));
 sky130_fd_sc_hd__a31oi_4 _24637_ (.A1(_00319_),
    .A2(_00321_),
    .A3(net210),
    .B1(_00323_),
    .Y(_00325_));
 sky130_fd_sc_hd__a21oi_1 _24638_ (.A1(_00322_),
    .A2(_00324_),
    .B1(net208),
    .Y(_00326_));
 sky130_fd_sc_hd__or3_1 _24639_ (.A(net231),
    .B(net228),
    .C(_00325_),
    .X(_00327_));
 sky130_fd_sc_hd__a31o_1 _24640_ (.A1(_00319_),
    .A2(_00321_),
    .A3(net210),
    .B1(net233),
    .X(_00329_));
 sky130_fd_sc_hd__a311oi_4 _24641_ (.A1(_00319_),
    .A2(_00321_),
    .A3(net210),
    .B1(_00323_),
    .C1(net233),
    .Y(_00330_));
 sky130_fd_sc_hd__nand3_1 _24642_ (.A(_00322_),
    .B(_00324_),
    .C(net235),
    .Y(_00331_));
 sky130_fd_sc_hd__a22oi_2 _24643_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_00322_),
    .B2(_00324_),
    .Y(_00332_));
 sky130_fd_sc_hd__a21o_2 _24644_ (.A1(_00322_),
    .A2(_00324_),
    .B1(net235),
    .X(_00333_));
 sky130_fd_sc_hd__o32a_1 _24645_ (.A1(net284),
    .A2(net282),
    .A3(_14410_),
    .B1(_14415_),
    .B2(_14419_),
    .X(_00334_));
 sky130_fd_sc_hd__a21oi_2 _24646_ (.A1(_14415_),
    .A2(_14418_),
    .B1(_14419_),
    .Y(_00335_));
 sky130_fd_sc_hd__o21a_2 _24647_ (.A1(_00330_),
    .A2(_00332_),
    .B1(_00335_),
    .X(_00336_));
 sky130_fd_sc_hd__o21ai_2 _24648_ (.A1(_00330_),
    .A2(_00332_),
    .B1(_00335_),
    .Y(_00337_));
 sky130_fd_sc_hd__o21ai_2 _24649_ (.A1(net235),
    .A2(_00325_),
    .B1(_00334_),
    .Y(_00338_));
 sky130_fd_sc_hd__o211ai_2 _24650_ (.A1(_00323_),
    .A2(_00329_),
    .B1(_00334_),
    .C1(_00333_),
    .Y(_00340_));
 sky130_fd_sc_hd__o22ai_4 _24651_ (.A1(net231),
    .A2(net228),
    .B1(_00330_),
    .B2(_00338_),
    .Y(_00341_));
 sky130_fd_sc_hd__o211ai_2 _24652_ (.A1(_00330_),
    .A2(_00338_),
    .B1(net208),
    .C1(_00337_),
    .Y(_00342_));
 sky130_fd_sc_hd__o22ai_4 _24653_ (.A1(net208),
    .A2(_00325_),
    .B1(_00336_),
    .B2(_00341_),
    .Y(_00343_));
 sky130_fd_sc_hd__o211a_1 _24654_ (.A1(net254),
    .A2(_14429_),
    .B1(_14055_),
    .C1(_14039_),
    .X(_00344_));
 sky130_fd_sc_hd__a21oi_1 _24655_ (.A1(_14039_),
    .A2(_14055_),
    .B1(_14434_),
    .Y(_00345_));
 sky130_fd_sc_hd__a31oi_2 _24656_ (.A1(_14039_),
    .A2(_14055_),
    .A3(_14433_),
    .B1(_14434_),
    .Y(_00346_));
 sky130_fd_sc_hd__a31oi_1 _24657_ (.A1(_00337_),
    .A2(_00340_),
    .A3(net208),
    .B1(net252),
    .Y(_00347_));
 sky130_fd_sc_hd__a311oi_4 _24658_ (.A1(_00337_),
    .A2(_00340_),
    .A3(net208),
    .B1(_00326_),
    .C1(net252),
    .Y(_00348_));
 sky130_fd_sc_hd__o221ai_4 _24659_ (.A1(net208),
    .A2(_00325_),
    .B1(_00336_),
    .B2(_00341_),
    .C1(_06314_),
    .Y(_00349_));
 sky130_fd_sc_hd__a2bb2oi_2 _24660_ (.A1_N(net284),
    .A2_N(net282),
    .B1(_00327_),
    .B2(_00342_),
    .Y(_00351_));
 sky130_fd_sc_hd__o21ai_2 _24661_ (.A1(net284),
    .A2(net282),
    .B1(_00343_),
    .Y(_00352_));
 sky130_fd_sc_hd__a21oi_1 _24662_ (.A1(_00327_),
    .A2(_00347_),
    .B1(_00351_),
    .Y(_00353_));
 sky130_fd_sc_hd__o211ai_2 _24663_ (.A1(_14434_),
    .A2(_00344_),
    .B1(_00349_),
    .C1(_00352_),
    .Y(_00354_));
 sky130_fd_sc_hd__o22ai_2 _24664_ (.A1(_14432_),
    .A2(_00345_),
    .B1(_00348_),
    .B2(_00351_),
    .Y(_00355_));
 sky130_fd_sc_hd__o211ai_4 _24665_ (.A1(net207),
    .A2(net206),
    .B1(_00354_),
    .C1(_00355_),
    .Y(_00356_));
 sky130_fd_sc_hd__a211o_2 _24666_ (.A1(_00327_),
    .A2(_00342_),
    .B1(net207),
    .C1(net205),
    .X(_00357_));
 sky130_fd_sc_hd__o211ai_2 _24667_ (.A1(_14432_),
    .A2(_00345_),
    .B1(_00349_),
    .C1(_00352_),
    .Y(_00358_));
 sky130_fd_sc_hd__o22ai_2 _24668_ (.A1(_14434_),
    .A2(_00344_),
    .B1(_00348_),
    .B2(_00351_),
    .Y(_00359_));
 sky130_fd_sc_hd__o211ai_4 _24669_ (.A1(net207),
    .A2(net205),
    .B1(_00358_),
    .C1(_00359_),
    .Y(_00360_));
 sky130_fd_sc_hd__nand2_1 _24670_ (.A(_00357_),
    .B(_00360_),
    .Y(_00362_));
 sky130_fd_sc_hd__o211a_1 _24671_ (.A1(_07233_),
    .A2(_00343_),
    .B1(_00356_),
    .C1(_06014_),
    .X(_00363_));
 sky130_fd_sc_hd__o211ai_4 _24672_ (.A1(_07233_),
    .A2(_00343_),
    .B1(_00356_),
    .C1(_06014_),
    .Y(_00364_));
 sky130_fd_sc_hd__and3_1 _24673_ (.A(_00360_),
    .B(net254),
    .C(_00357_),
    .X(_00365_));
 sky130_fd_sc_hd__o211ai_4 _24674_ (.A1(net285),
    .A2(_06012_),
    .B1(_00357_),
    .C1(_00360_),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2_1 _24675_ (.A(_00364_),
    .B(_00366_),
    .Y(_00367_));
 sky130_fd_sc_hd__a22oi_2 _24676_ (.A1(_05768_),
    .A2(_14446_),
    .B1(_14460_),
    .B2(_14462_),
    .Y(_00368_));
 sky130_fd_sc_hd__o22ai_4 _24677_ (.A1(net263),
    .A2(_14448_),
    .B1(_00002_),
    .B2(_14459_),
    .Y(_00369_));
 sky130_fd_sc_hd__o21ai_4 _24678_ (.A1(_14452_),
    .A2(_00368_),
    .B1(_00367_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand3_4 _24679_ (.A(_00369_),
    .B(_00366_),
    .C(_00364_),
    .Y(_00371_));
 sky130_fd_sc_hd__nand3_1 _24680_ (.A(_00370_),
    .B(_00371_),
    .C(net163),
    .Y(_00373_));
 sky130_fd_sc_hd__o311a_4 _24681_ (.A1(net207),
    .A2(_00343_),
    .A3(net206),
    .B1(_07550_),
    .C1(_00356_),
    .X(_00374_));
 sky130_fd_sc_hd__a211o_1 _24682_ (.A1(_00357_),
    .A2(_00360_),
    .B1(_07544_),
    .C1(_07546_),
    .X(_00375_));
 sky130_fd_sc_hd__a31oi_2 _24683_ (.A1(_00370_),
    .A2(_00371_),
    .A3(net163),
    .B1(_00374_),
    .Y(_00376_));
 sky130_fd_sc_hd__a311o_1 _24684_ (.A1(_00370_),
    .A2(_00371_),
    .A3(net163),
    .B1(_00374_),
    .C1(net161),
    .X(_00377_));
 sky130_fd_sc_hd__a22oi_2 _24685_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_00373_),
    .B2(_00375_),
    .Y(_00378_));
 sky130_fd_sc_hd__a22o_1 _24686_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_00373_),
    .B2(_00375_),
    .X(_00379_));
 sky130_fd_sc_hd__a31o_1 _24687_ (.A1(_00370_),
    .A2(_00371_),
    .A3(net163),
    .B1(_05768_),
    .X(_00380_));
 sky130_fd_sc_hd__a311oi_4 _24688_ (.A1(_00370_),
    .A2(_00371_),
    .A3(net163),
    .B1(_00374_),
    .C1(_05768_),
    .Y(_00381_));
 sky130_fd_sc_hd__a311o_1 _24689_ (.A1(_00370_),
    .A2(_00371_),
    .A3(net163),
    .B1(_00374_),
    .C1(_05768_),
    .X(_00382_));
 sky130_fd_sc_hd__o21ai_1 _24690_ (.A1(_14082_),
    .A2(_00014_),
    .B1(_00013_),
    .Y(_00384_));
 sky130_fd_sc_hd__a21boi_2 _24691_ (.A1(_00013_),
    .A2(_00017_),
    .B1_N(_00012_),
    .Y(_00385_));
 sky130_fd_sc_hd__o2bb2ai_4 _24692_ (.A1_N(_00013_),
    .A2_N(_00017_),
    .B1(_14467_),
    .B2(_00010_),
    .Y(_00386_));
 sky130_fd_sc_hd__o211ai_1 _24693_ (.A1(_00374_),
    .A2(_00380_),
    .B1(_00386_),
    .C1(_00379_),
    .Y(_00387_));
 sky130_fd_sc_hd__o21ai_1 _24694_ (.A1(_00378_),
    .A2(_00381_),
    .B1(_00385_),
    .Y(_00388_));
 sky130_fd_sc_hd__o211ai_2 _24695_ (.A1(net183),
    .A2(net182),
    .B1(_00387_),
    .C1(_00388_),
    .Y(_00389_));
 sky130_fd_sc_hd__a21oi_1 _24696_ (.A1(_00373_),
    .A2(_00375_),
    .B1(net161),
    .Y(_00390_));
 sky130_fd_sc_hd__or3_2 _24697_ (.A(net183),
    .B(net182),
    .C(_00376_),
    .X(_00391_));
 sky130_fd_sc_hd__o21ai_2 _24698_ (.A1(_00378_),
    .A2(_00381_),
    .B1(_00386_),
    .Y(_00392_));
 sky130_fd_sc_hd__o211ai_4 _24699_ (.A1(_00374_),
    .A2(_00380_),
    .B1(_00385_),
    .C1(_00379_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand3_2 _24700_ (.A(_00392_),
    .B(_00393_),
    .C(net161),
    .Y(_00395_));
 sky130_fd_sc_hd__and3_2 _24701_ (.A(_08301_),
    .B(_00377_),
    .C(_00389_),
    .X(_00396_));
 sky130_fd_sc_hd__a211o_1 _24702_ (.A1(_00391_),
    .A2(_00395_),
    .B1(_08296_),
    .C1(net179),
    .X(_00397_));
 sky130_fd_sc_hd__a311oi_4 _24703_ (.A1(_00392_),
    .A2(_00393_),
    .A3(net161),
    .B1(_00390_),
    .C1(net292),
    .Y(_00398_));
 sky130_fd_sc_hd__nand3_4 _24704_ (.A(_00395_),
    .B(_05507_),
    .C(_00391_),
    .Y(_00399_));
 sky130_fd_sc_hd__o211ai_4 _24705_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_00377_),
    .C1(_00389_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2_1 _24706_ (.A(_00399_),
    .B(_00400_),
    .Y(_00401_));
 sky130_fd_sc_hd__a21oi_1 _24707_ (.A1(net294),
    .A2(_00026_),
    .B1(_00030_),
    .Y(_00402_));
 sky130_fd_sc_hd__o21ai_1 _24708_ (.A1(_00031_),
    .A2(_00032_),
    .B1(_00036_),
    .Y(_00403_));
 sky130_fd_sc_hd__a21oi_2 _24709_ (.A1(_00034_),
    .A2(_00030_),
    .B1(_00035_),
    .Y(_00404_));
 sky130_fd_sc_hd__o2bb2ai_4 _24710_ (.A1_N(_00399_),
    .A2_N(_00400_),
    .B1(_00402_),
    .B2(_00032_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand3_4 _24711_ (.A(_00403_),
    .B(_00400_),
    .C(_00399_),
    .Y(_00407_));
 sky130_fd_sc_hd__nand3_1 _24712_ (.A(_00406_),
    .B(_00407_),
    .C(net159),
    .Y(_00408_));
 sky130_fd_sc_hd__a31oi_4 _24713_ (.A1(_00406_),
    .A2(_00407_),
    .A3(net159),
    .B1(_00396_),
    .Y(_00409_));
 sky130_fd_sc_hd__a31o_1 _24714_ (.A1(_00406_),
    .A2(_00407_),
    .A3(net159),
    .B1(_00396_),
    .X(_00410_));
 sky130_fd_sc_hd__a31oi_2 _24715_ (.A1(_04238_),
    .A2(_00027_),
    .A3(_00039_),
    .B1(_00051_),
    .Y(_00411_));
 sky130_fd_sc_hd__a31o_1 _24716_ (.A1(_04227_),
    .A2(_00041_),
    .A3(_00045_),
    .B1(_00052_),
    .X(_00412_));
 sky130_fd_sc_hd__a32oi_2 _24717_ (.A1(_04227_),
    .A2(_00041_),
    .A3(_00045_),
    .B1(_00047_),
    .B2(_00052_),
    .Y(_00413_));
 sky130_fd_sc_hd__a31o_1 _24718_ (.A1(_00406_),
    .A2(_00407_),
    .A3(net159),
    .B1(_05249_),
    .X(_00414_));
 sky130_fd_sc_hd__a311oi_4 _24719_ (.A1(_00406_),
    .A2(_00407_),
    .A3(net159),
    .B1(_00396_),
    .C1(net294),
    .Y(_00415_));
 sky130_fd_sc_hd__a2bb2oi_2 _24720_ (.A1_N(net318),
    .A2_N(net315),
    .B1(_00397_),
    .B2(_00408_),
    .Y(_00417_));
 sky130_fd_sc_hd__a22o_1 _24721_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_00397_),
    .B2(_00408_),
    .X(_00418_));
 sky130_fd_sc_hd__o221ai_1 _24722_ (.A1(_00048_),
    .A2(_00411_),
    .B1(_00414_),
    .B2(_00396_),
    .C1(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__o2bb2ai_1 _24723_ (.A1_N(_00047_),
    .A2_N(_00412_),
    .B1(_00415_),
    .B2(_00417_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand3_1 _24724_ (.A(_00419_),
    .B(_00420_),
    .C(net149),
    .Y(_00421_));
 sky130_fd_sc_hd__or3_1 _24725_ (.A(net158),
    .B(_08712_),
    .C(_00409_),
    .X(_00422_));
 sky130_fd_sc_hd__o21ai_1 _24726_ (.A1(net295),
    .A2(_00409_),
    .B1(_00413_),
    .Y(_00423_));
 sky130_fd_sc_hd__o22ai_2 _24727_ (.A1(_00048_),
    .A2(_00411_),
    .B1(_00415_),
    .B2(_00417_),
    .Y(_00424_));
 sky130_fd_sc_hd__o221ai_4 _24728_ (.A1(net158),
    .A2(_08712_),
    .B1(_00415_),
    .B2(_00423_),
    .C1(_00424_),
    .Y(_00425_));
 sky130_fd_sc_hd__o21ai_2 _24729_ (.A1(_08714_),
    .A2(_00409_),
    .B1(_00425_),
    .Y(_00426_));
 sky130_fd_sc_hd__a2bb2oi_1 _24730_ (.A1_N(net340),
    .A2_N(_04184_),
    .B1(_00422_),
    .B2(_00425_),
    .Y(_00428_));
 sky130_fd_sc_hd__o211ai_4 _24731_ (.A1(_00410_),
    .A2(net149),
    .B1(_04238_),
    .C1(_00421_),
    .Y(_00429_));
 sky130_fd_sc_hd__o211a_1 _24732_ (.A1(_08714_),
    .A2(_00409_),
    .B1(_04227_),
    .C1(_00425_),
    .X(_00430_));
 sky130_fd_sc_hd__o211ai_4 _24733_ (.A1(_08714_),
    .A2(_00409_),
    .B1(_04227_),
    .C1(_00425_),
    .Y(_00431_));
 sky130_fd_sc_hd__a21oi_1 _24734_ (.A1(_00068_),
    .A2(_00071_),
    .B1(_00061_),
    .Y(_00432_));
 sky130_fd_sc_hd__a32o_1 _24735_ (.A1(_02104_),
    .A2(_02126_),
    .A3(_00060_),
    .B1(_00068_),
    .B2(_00071_),
    .X(_00433_));
 sky130_fd_sc_hd__o2111ai_4 _24736_ (.A1(_00063_),
    .A2(_00073_),
    .B1(_00429_),
    .C1(_00431_),
    .D1(_00062_),
    .Y(_00434_));
 sky130_fd_sc_hd__o2bb2ai_1 _24737_ (.A1_N(_00062_),
    .A2_N(_00075_),
    .B1(_00428_),
    .B2(_00430_),
    .Y(_00435_));
 sky130_fd_sc_hd__o211ai_4 _24738_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_00434_),
    .C1(_00435_),
    .Y(_00436_));
 sky130_fd_sc_hd__a211o_1 _24739_ (.A1(_00422_),
    .A2(_00425_),
    .B1(_09120_),
    .C1(_09121_),
    .X(_00437_));
 sky130_fd_sc_hd__o2bb2ai_1 _24740_ (.A1_N(_00429_),
    .A2_N(_00431_),
    .B1(_00432_),
    .B2(_00063_),
    .Y(_00439_));
 sky130_fd_sc_hd__o2111ai_1 _24741_ (.A1(_02148_),
    .A2(_00060_),
    .B1(_00429_),
    .C1(_00431_),
    .D1(_00433_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand3_1 _24742_ (.A(_09125_),
    .B(_00439_),
    .C(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__o21ai_4 _24743_ (.A1(net146),
    .A2(_00426_),
    .B1(_00436_),
    .Y(_00442_));
 sky130_fd_sc_hd__o21ai_2 _24744_ (.A1(_09559_),
    .A2(_09560_),
    .B1(_00442_),
    .Y(_00443_));
 sky130_fd_sc_hd__o211a_2 _24745_ (.A1(_00426_),
    .A2(_09125_),
    .B1(_02148_),
    .C1(_00436_),
    .X(_00444_));
 sky130_fd_sc_hd__o211ai_1 _24746_ (.A1(_00426_),
    .A2(net146),
    .B1(_02148_),
    .C1(_00436_),
    .Y(_00445_));
 sky130_fd_sc_hd__and3_1 _24747_ (.A(_00441_),
    .B(_02137_),
    .C(_00437_),
    .X(_00446_));
 sky130_fd_sc_hd__nand3_2 _24748_ (.A(_00441_),
    .B(_02137_),
    .C(_00437_),
    .Y(_00447_));
 sky130_fd_sc_hd__nand2_1 _24749_ (.A(_00445_),
    .B(_00447_),
    .Y(_00448_));
 sky130_fd_sc_hd__a211oi_1 _24750_ (.A1(_13726_),
    .A2(_13716_),
    .B1(_13289_),
    .C1(_13724_),
    .Y(_00450_));
 sky130_fd_sc_hd__o211ai_2 _24751_ (.A1(_14126_),
    .A2(_14149_),
    .B1(_00450_),
    .C1(_14153_),
    .Y(_00451_));
 sky130_fd_sc_hd__a31oi_4 _24752_ (.A1(_00078_),
    .A2(_00080_),
    .A3(_00240_),
    .B1(_00451_),
    .Y(_00452_));
 sky130_fd_sc_hd__a31o_1 _24753_ (.A1(_00078_),
    .A2(_00080_),
    .A3(_00240_),
    .B1(_00451_),
    .X(_00453_));
 sky130_fd_sc_hd__a211oi_1 _24754_ (.A1(_00089_),
    .A2(_00085_),
    .B1(_00086_),
    .C1(_00452_),
    .Y(_00454_));
 sky130_fd_sc_hd__o211ai_4 _24755_ (.A1(_00090_),
    .A2(_00084_),
    .B1(_00087_),
    .C1(_00453_),
    .Y(_00455_));
 sky130_fd_sc_hd__o211a_1 _24756_ (.A1(_00240_),
    .A2(_00081_),
    .B1(_00452_),
    .C1(_13291_),
    .X(_00456_));
 sky130_fd_sc_hd__o211ai_4 _24757_ (.A1(_00240_),
    .A2(_00081_),
    .B1(_00452_),
    .C1(_13291_),
    .Y(_00457_));
 sky130_fd_sc_hd__nor2_1 _24758_ (.A(_00454_),
    .B(_00456_),
    .Y(_00458_));
 sky130_fd_sc_hd__inv_2 _24759_ (.A(_00458_),
    .Y(_00459_));
 sky130_fd_sc_hd__nand3_2 _24760_ (.A(_00447_),
    .B(_00455_),
    .C(_00457_),
    .Y(_00461_));
 sky130_fd_sc_hd__o22ai_2 _24761_ (.A1(_00444_),
    .A2(_00446_),
    .B1(_00454_),
    .B2(_00456_),
    .Y(_00462_));
 sky130_fd_sc_hd__a21o_1 _24762_ (.A1(_00455_),
    .A2(_00457_),
    .B1(_00448_),
    .X(_00463_));
 sky130_fd_sc_hd__o211ai_1 _24763_ (.A1(_00444_),
    .A2(_00446_),
    .B1(_00455_),
    .C1(_00457_),
    .Y(_00464_));
 sky130_fd_sc_hd__nand3_1 _24764_ (.A(net143),
    .B(_00463_),
    .C(_00464_),
    .Y(_00465_));
 sky130_fd_sc_hd__or3_1 _24765_ (.A(_09553_),
    .B(net155),
    .C(_00442_),
    .X(_00466_));
 sky130_fd_sc_hd__o221ai_4 _24766_ (.A1(_09553_),
    .A2(net155),
    .B1(_00444_),
    .B2(_00461_),
    .C1(_00462_),
    .Y(_00467_));
 sky130_fd_sc_hd__and3_1 _24767_ (.A(_00465_),
    .B(_09578_),
    .C(_00443_),
    .X(_00468_));
 sky130_fd_sc_hd__a22o_1 _24768_ (.A1(_09575_),
    .A2(_09577_),
    .B1(_00466_),
    .B2(_00467_),
    .X(_00469_));
 sky130_fd_sc_hd__o311a_1 _24769_ (.A1(_09553_),
    .A2(net155),
    .A3(_00442_),
    .B1(_00240_),
    .C1(_00467_),
    .X(_00470_));
 sky130_fd_sc_hd__o211ai_4 _24770_ (.A1(net143),
    .A2(_00442_),
    .B1(_00240_),
    .C1(_00467_),
    .Y(_00472_));
 sky130_fd_sc_hd__a2bb2oi_1 _24771_ (.A1_N(_00174_),
    .A2_N(net344),
    .B1(_00466_),
    .B2(_00467_),
    .Y(_00473_));
 sky130_fd_sc_hd__o211ai_4 _24772_ (.A1(_00174_),
    .A2(net344),
    .B1(_00443_),
    .C1(_00465_),
    .Y(_00474_));
 sky130_fd_sc_hd__o221a_1 _24773_ (.A1(_14166_),
    .A2(_14163_),
    .B1(_12888_),
    .B2(_00094_),
    .C1(_14161_),
    .X(_00475_));
 sky130_fd_sc_hd__o32a_1 _24774_ (.A1(net361),
    .A2(net345),
    .A3(_00095_),
    .B1(_00098_),
    .B2(_00101_),
    .X(_00476_));
 sky130_fd_sc_hd__a21oi_2 _24775_ (.A1(_00098_),
    .A2(_00100_),
    .B1(_00101_),
    .Y(_00477_));
 sky130_fd_sc_hd__o2bb2ai_2 _24776_ (.A1_N(_00472_),
    .A2_N(_00474_),
    .B1(_00475_),
    .B2(_00099_),
    .Y(_00478_));
 sky130_fd_sc_hd__nand3_1 _24777_ (.A(_00476_),
    .B(_00474_),
    .C(_00472_),
    .Y(_00479_));
 sky130_fd_sc_hd__o311a_1 _24778_ (.A1(_00477_),
    .A2(_00473_),
    .A3(_00470_),
    .B1(_09579_),
    .C1(_00478_),
    .X(_00480_));
 sky130_fd_sc_hd__nand3_2 _24779_ (.A(_09579_),
    .B(_00478_),
    .C(_00479_),
    .Y(_00481_));
 sky130_fd_sc_hd__o311a_1 _24780_ (.A1(net365),
    .A2(net362),
    .A3(_14172_),
    .B1(_14185_),
    .C1(_00112_),
    .X(_00483_));
 sky130_fd_sc_hd__a31oi_2 _24781_ (.A1(_14175_),
    .A2(_14185_),
    .A3(_00112_),
    .B1(_00113_),
    .Y(_00484_));
 sky130_fd_sc_hd__a311oi_2 _24782_ (.A1(_09579_),
    .A2(_00478_),
    .A3(_00479_),
    .B1(_00468_),
    .C1(_12899_),
    .Y(_00485_));
 sky130_fd_sc_hd__o211ai_2 _24783_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_00469_),
    .C1(_00481_),
    .Y(_00486_));
 sky130_fd_sc_hd__a21oi_2 _24784_ (.A1(_00469_),
    .A2(_00481_),
    .B1(_12888_),
    .Y(_00487_));
 sky130_fd_sc_hd__o21ai_1 _24785_ (.A1(_00468_),
    .A2(_00480_),
    .B1(_12899_),
    .Y(_00488_));
 sky130_fd_sc_hd__nand3_1 _24786_ (.A(_00488_),
    .B(_00484_),
    .C(_00486_),
    .Y(_00489_));
 sky130_fd_sc_hd__o22ai_1 _24787_ (.A1(_00113_),
    .A2(_00483_),
    .B1(_00485_),
    .B2(_00487_),
    .Y(_00490_));
 sky130_fd_sc_hd__a211o_1 _24788_ (.A1(_00469_),
    .A2(_00481_),
    .B1(_10474_),
    .C1(net138),
    .X(_00491_));
 sky130_fd_sc_hd__o211ai_2 _24789_ (.A1(_10474_),
    .A2(net138),
    .B1(_00489_),
    .C1(_00490_),
    .Y(_00492_));
 sky130_fd_sc_hd__o21ai_1 _24790_ (.A1(_00124_),
    .A2(_00122_),
    .B1(_00121_),
    .Y(_00494_));
 sky130_fd_sc_hd__and3_1 _24791_ (.A(_00492_),
    .B(_11298_),
    .C(_00491_),
    .X(_00495_));
 sky130_fd_sc_hd__o211ai_1 _24792_ (.A1(_11254_),
    .A2(_11276_),
    .B1(_00491_),
    .C1(_00492_),
    .Y(_00496_));
 sky130_fd_sc_hd__a21oi_1 _24793_ (.A1(_00491_),
    .A2(_00492_),
    .B1(_11298_),
    .Y(_00497_));
 sky130_fd_sc_hd__a22o_1 _24794_ (.A1(_11221_),
    .A2(_11243_),
    .B1(_00491_),
    .B2(_00492_),
    .X(_00498_));
 sky130_fd_sc_hd__a211o_1 _24795_ (.A1(_00491_),
    .A2(_00492_),
    .B1(_10949_),
    .C1(net136),
    .X(_00499_));
 sky130_fd_sc_hd__nand2_1 _24796_ (.A(_00498_),
    .B(_00494_),
    .Y(_00500_));
 sky130_fd_sc_hd__o221ai_2 _24797_ (.A1(_00124_),
    .A2(_00122_),
    .B1(_00497_),
    .B2(_00495_),
    .C1(_00121_),
    .Y(_00501_));
 sky130_fd_sc_hd__o211ai_2 _24798_ (.A1(_00495_),
    .A2(_00500_),
    .B1(_00501_),
    .C1(_10954_),
    .Y(_00502_));
 sky130_fd_sc_hd__nand4_2 _24799_ (.A(_11460_),
    .B(_11462_),
    .C(_00499_),
    .D(_00502_),
    .Y(_00503_));
 sky130_fd_sc_hd__a21oi_1 _24800_ (.A1(_00499_),
    .A2(_00502_),
    .B1(_10015_),
    .Y(_00505_));
 sky130_fd_sc_hd__o211ai_2 _24801_ (.A1(net365),
    .A2(net362),
    .B1(_00499_),
    .C1(_00502_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2b_1 _24802_ (.A_N(_00505_),
    .B(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__o21ai_2 _24803_ (.A1(_00128_),
    .A2(_00129_),
    .B1(_00132_),
    .Y(_00508_));
 sky130_fd_sc_hd__a21oi_1 _24804_ (.A1(_00507_),
    .A2(_00508_),
    .B1(_11464_),
    .Y(_00509_));
 sky130_fd_sc_hd__o21ai_1 _24805_ (.A1(_00507_),
    .A2(_00508_),
    .B1(_00509_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _24806_ (.A(_00503_),
    .B(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__and3_1 _24807_ (.A(_08918_),
    .B(_00503_),
    .C(_00510_),
    .X(_00512_));
 sky130_fd_sc_hd__a21o_1 _24808_ (.A1(_00503_),
    .A2(_00510_),
    .B1(_08918_),
    .X(_00513_));
 sky130_fd_sc_hd__and2b_1 _24809_ (.A_N(_00512_),
    .B(_00513_),
    .X(_00514_));
 sky130_fd_sc_hd__a21o_1 _24810_ (.A1(_00136_),
    .A2(_00137_),
    .B1(_00138_),
    .X(_00516_));
 sky130_fd_sc_hd__or2_1 _24811_ (.A(_00516_),
    .B(_00514_),
    .X(_00517_));
 sky130_fd_sc_hd__a21bo_1 _24812_ (.A1(_00517_),
    .A2(_11943_),
    .B1_N(_00511_),
    .X(_00518_));
 sky130_fd_sc_hd__a21oi_1 _24813_ (.A1(_05119_),
    .A2(_00145_),
    .B1(_00518_),
    .Y(_00519_));
 sky130_fd_sc_hd__and3_1 _24814_ (.A(_05119_),
    .B(_00145_),
    .C(_00518_),
    .X(_00520_));
 sky130_fd_sc_hd__nor2_1 _24815_ (.A(_00519_),
    .B(_00520_),
    .Y(net96));
 sky130_fd_sc_hd__or2_1 _24816_ (.A(_00145_),
    .B(_00518_),
    .X(_00521_));
 sky130_fd_sc_hd__o311a_1 _24817_ (.A1(_03399_),
    .A2(net24),
    .A3(_10962_),
    .B1(_00149_),
    .C1(_00155_),
    .X(_00522_));
 sky130_fd_sc_hd__a31o_1 _24818_ (.A1(_11471_),
    .A2(_00149_),
    .A3(_00155_),
    .B1(_11079_),
    .X(_00523_));
 sky130_fd_sc_hd__or4_1 _24819_ (.A(_11079_),
    .B(net329),
    .C(net327),
    .D(_00522_),
    .X(_00524_));
 sky130_fd_sc_hd__a311o_1 _24820_ (.A1(_11471_),
    .A2(_00149_),
    .A3(_00155_),
    .B1(_10970_),
    .C1(_11079_),
    .X(_00526_));
 sky130_fd_sc_hd__o21ai_1 _24821_ (.A1(_11079_),
    .A2(_00522_),
    .B1(_10970_),
    .Y(_00527_));
 sky130_fd_sc_hd__and2_1 _24822_ (.A(_00526_),
    .B(_00527_),
    .X(_00528_));
 sky130_fd_sc_hd__nand2_1 _24823_ (.A(_00526_),
    .B(_00527_),
    .Y(_00529_));
 sky130_fd_sc_hd__o21ai_1 _24824_ (.A1(_00162_),
    .A2(_00165_),
    .B1(_00160_),
    .Y(_00530_));
 sky130_fd_sc_hd__a21oi_2 _24825_ (.A1(_00160_),
    .A2(_00168_),
    .B1(_00529_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _24826_ (.A(_00530_),
    .B(_00528_),
    .Y(_00532_));
 sky130_fd_sc_hd__o211ai_1 _24827_ (.A1(_00162_),
    .A2(_00165_),
    .B1(_00529_),
    .C1(_00160_),
    .Y(_00533_));
 sky130_fd_sc_hd__o21ai_2 _24828_ (.A1(net329),
    .A2(net327),
    .B1(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__o221ai_1 _24829_ (.A1(net329),
    .A2(net327),
    .B1(_00528_),
    .B2(_00530_),
    .C1(_00532_),
    .Y(_00535_));
 sky130_fd_sc_hd__o32a_2 _24830_ (.A1(_11079_),
    .A2(net311),
    .A3(_00522_),
    .B1(_00534_),
    .B2(_00531_),
    .X(_00537_));
 sky130_fd_sc_hd__o22ai_1 _24831_ (.A1(net311),
    .A2(_00523_),
    .B1(_00534_),
    .B2(_00531_),
    .Y(_00538_));
 sky130_fd_sc_hd__a2bb2oi_1 _24832_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_00524_),
    .B2(_00535_),
    .Y(_00539_));
 sky130_fd_sc_hd__o21ai_2 _24833_ (.A1(_10487_),
    .A2(net166),
    .B1(_00538_),
    .Y(_00540_));
 sky130_fd_sc_hd__o221a_1 _24834_ (.A1(net311),
    .A2(_00523_),
    .B1(_00534_),
    .B2(_00531_),
    .C1(net150),
    .X(_00541_));
 sky130_fd_sc_hd__o221ai_1 _24835_ (.A1(net311),
    .A2(_00523_),
    .B1(_00534_),
    .B2(_00531_),
    .C1(net150),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_1 _24836_ (.A(_00540_),
    .B(_00542_),
    .Y(_00543_));
 sky130_fd_sc_hd__a31oi_4 _24837_ (.A1(_00177_),
    .A2(_00181_),
    .A3(_00183_),
    .B1(_00175_),
    .Y(_00544_));
 sky130_fd_sc_hd__o221a_2 _24838_ (.A1(net153),
    .A2(_00171_),
    .B1(_00539_),
    .B2(_00541_),
    .C1(_00188_),
    .X(_00545_));
 sky130_fd_sc_hd__o22ai_4 _24839_ (.A1(_00011_),
    .A2(net321),
    .B1(_00544_),
    .B2(_00543_),
    .Y(_00546_));
 sky130_fd_sc_hd__o22ai_4 _24840_ (.A1(net307),
    .A2(_00537_),
    .B1(_00545_),
    .B2(_00546_),
    .Y(_00548_));
 sky130_fd_sc_hd__o21a_1 _24841_ (.A1(_01919_),
    .A2(_01930_),
    .B1(_00548_),
    .X(_00549_));
 sky130_fd_sc_hd__o21ai_2 _24842_ (.A1(_01919_),
    .A2(_01930_),
    .B1(_00548_),
    .Y(_00550_));
 sky130_fd_sc_hd__o221ai_4 _24843_ (.A1(net307),
    .A2(_00537_),
    .B1(_00545_),
    .B2(_00546_),
    .C1(net153),
    .Y(_00551_));
 sky130_fd_sc_hd__o21a_1 _24844_ (.A1(net170),
    .A2(net169),
    .B1(_00548_),
    .X(_00552_));
 sky130_fd_sc_hd__o21ai_2 _24845_ (.A1(net170),
    .A2(net169),
    .B1(_00548_),
    .Y(_00553_));
 sky130_fd_sc_hd__and3_1 _24846_ (.A(_13432_),
    .B(_13870_),
    .C(_13871_),
    .X(_00554_));
 sky130_fd_sc_hd__nand3_1 _24847_ (.A(_00195_),
    .B(_00554_),
    .C(_14275_),
    .Y(_00555_));
 sky130_fd_sc_hd__o211ai_4 _24848_ (.A1(_00200_),
    .A2(_00194_),
    .B1(_00198_),
    .C1(_00555_),
    .Y(_00556_));
 sky130_fd_sc_hd__nand4_1 _24849_ (.A(_00554_),
    .B(_14274_),
    .C(_14272_),
    .D(_13443_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand3b_4 _24850_ (.A_N(_00557_),
    .B(_00198_),
    .C(_00195_),
    .Y(_00559_));
 sky130_fd_sc_hd__a22oi_1 _24851_ (.A1(_00551_),
    .A2(_00553_),
    .B1(_00556_),
    .B2(_00559_),
    .Y(_00560_));
 sky130_fd_sc_hd__a22o_1 _24852_ (.A1(_00551_),
    .A2(_00553_),
    .B1(_00556_),
    .B2(_00559_),
    .X(_00561_));
 sky130_fd_sc_hd__and4_1 _24853_ (.A(_00551_),
    .B(_00553_),
    .C(_00556_),
    .D(_00559_),
    .X(_00562_));
 sky130_fd_sc_hd__nand4_2 _24854_ (.A(_00551_),
    .B(_00553_),
    .C(_00556_),
    .D(_00559_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand3_2 _24855_ (.A(_00561_),
    .B(_00563_),
    .C(net278),
    .Y(_00564_));
 sky130_fd_sc_hd__o22ai_2 _24856_ (.A1(net304),
    .A2(_01951_),
    .B1(_00560_),
    .B2(_00562_),
    .Y(_00565_));
 sky130_fd_sc_hd__o311a_2 _24857_ (.A1(net304),
    .A2(_00548_),
    .A3(_01951_),
    .B1(_04040_),
    .C1(_00565_),
    .X(_00566_));
 sky130_fd_sc_hd__a211o_2 _24858_ (.A1(_00550_),
    .A2(_00564_),
    .B1(net302),
    .C1(_04019_),
    .X(_00567_));
 sky130_fd_sc_hd__a311oi_4 _24859_ (.A1(_00561_),
    .A2(_00563_),
    .A3(net278),
    .B1(_09595_),
    .C1(_00549_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand3_2 _24860_ (.A(_00564_),
    .B(net172),
    .C(_00550_),
    .Y(_00570_));
 sky130_fd_sc_hd__a22oi_2 _24861_ (.A1(_09589_),
    .A2(_09591_),
    .B1(_00550_),
    .B2(_00564_),
    .Y(_00571_));
 sky130_fd_sc_hd__o211ai_4 _24862_ (.A1(_00548_),
    .A2(net278),
    .B1(_09595_),
    .C1(_00565_),
    .Y(_00572_));
 sky130_fd_sc_hd__o32a_1 _24863_ (.A1(_09134_),
    .A2(_09135_),
    .A3(_00205_),
    .B1(_00211_),
    .B2(_00208_),
    .X(_00573_));
 sky130_fd_sc_hd__o32ai_4 _24864_ (.A1(_09134_),
    .A2(_09135_),
    .A3(_00205_),
    .B1(_00211_),
    .B2(_00208_),
    .Y(_00574_));
 sky130_fd_sc_hd__o21ai_4 _24865_ (.A1(_00568_),
    .A2(_00571_),
    .B1(_00574_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand3_2 _24866_ (.A(_00573_),
    .B(_00572_),
    .C(_00570_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand3_2 _24867_ (.A(_00575_),
    .B(_00576_),
    .C(_04029_),
    .Y(_00577_));
 sky130_fd_sc_hd__a31o_2 _24868_ (.A1(_00575_),
    .A2(_00576_),
    .A3(_04029_),
    .B1(_00566_),
    .X(_00578_));
 sky130_fd_sc_hd__o221a_1 _24869_ (.A1(net199),
    .A2(_14301_),
    .B1(net177),
    .B2(_00220_),
    .C1(_00226_),
    .X(_00579_));
 sky130_fd_sc_hd__o21ai_1 _24870_ (.A1(net177),
    .A2(_00220_),
    .B1(_00228_),
    .Y(_00581_));
 sky130_fd_sc_hd__a22oi_1 _24871_ (.A1(net177),
    .A2(_00220_),
    .B1(_00226_),
    .B2(_14313_),
    .Y(_00582_));
 sky130_fd_sc_hd__o21ai_1 _24872_ (.A1(_00223_),
    .A2(_00228_),
    .B1(_00222_),
    .Y(_00583_));
 sky130_fd_sc_hd__a31o_1 _24873_ (.A1(_00575_),
    .A2(_00576_),
    .A3(_04029_),
    .B1(net173),
    .X(_00584_));
 sky130_fd_sc_hd__a311oi_4 _24874_ (.A1(_00575_),
    .A2(_00576_),
    .A3(_04029_),
    .B1(net173),
    .C1(_00566_),
    .Y(_00585_));
 sky130_fd_sc_hd__o211ai_2 _24875_ (.A1(_09136_),
    .A2(_09138_),
    .B1(_00567_),
    .C1(_00577_),
    .Y(_00586_));
 sky130_fd_sc_hd__a2bb2oi_4 _24876_ (.A1_N(_09134_),
    .A2_N(net192),
    .B1(_00567_),
    .B2(_00577_),
    .Y(_00587_));
 sky130_fd_sc_hd__a2bb2o_1 _24877_ (.A1_N(_09134_),
    .A2_N(net192),
    .B1(_00567_),
    .B2(_00577_),
    .X(_00588_));
 sky130_fd_sc_hd__nor2_1 _24878_ (.A(_00585_),
    .B(_00587_),
    .Y(_00589_));
 sky130_fd_sc_hd__o211ai_1 _24879_ (.A1(_00223_),
    .A2(_00579_),
    .B1(_00586_),
    .C1(_00588_),
    .Y(_00590_));
 sky130_fd_sc_hd__o22ai_1 _24880_ (.A1(_00221_),
    .A2(_00582_),
    .B1(_00585_),
    .B2(_00587_),
    .Y(_00592_));
 sky130_fd_sc_hd__nand3_2 _24881_ (.A(_00590_),
    .B(_00592_),
    .C(net271),
    .Y(_00593_));
 sky130_fd_sc_hd__a211o_1 _24882_ (.A1(_00567_),
    .A2(_00577_),
    .B1(net296),
    .C1(_05232_),
    .X(_00594_));
 sky130_fd_sc_hd__o211ai_1 _24883_ (.A1(_00221_),
    .A2(_00582_),
    .B1(_00586_),
    .C1(_00588_),
    .Y(_00595_));
 sky130_fd_sc_hd__o22ai_1 _24884_ (.A1(_00223_),
    .A2(_00579_),
    .B1(_00585_),
    .B2(_00587_),
    .Y(_00596_));
 sky130_fd_sc_hd__nand3_2 _24885_ (.A(_00595_),
    .B(_00596_),
    .C(net271),
    .Y(_00597_));
 sky130_fd_sc_hd__o21ai_2 _24886_ (.A1(net271),
    .A2(_00578_),
    .B1(_00593_),
    .Y(_00598_));
 sky130_fd_sc_hd__inv_2 _24887_ (.A(_00598_),
    .Y(_00599_));
 sky130_fd_sc_hd__and3_2 _24888_ (.A(_05486_),
    .B(_00594_),
    .C(_00597_),
    .X(_00600_));
 sky130_fd_sc_hd__o211a_1 _24889_ (.A1(_00578_),
    .A2(net271),
    .B1(net175),
    .C1(_00593_),
    .X(_00601_));
 sky130_fd_sc_hd__o211ai_4 _24890_ (.A1(_00578_),
    .A2(net271),
    .B1(net175),
    .C1(_00593_),
    .Y(_00603_));
 sky130_fd_sc_hd__and3_1 _24891_ (.A(_00597_),
    .B(net177),
    .C(_00594_),
    .X(_00604_));
 sky130_fd_sc_hd__nand3_4 _24892_ (.A(_00597_),
    .B(net177),
    .C(_00594_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_1 _24893_ (.A(_00603_),
    .B(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__a22oi_2 _24894_ (.A1(net198),
    .A2(_00236_),
    .B1(_00249_),
    .B2(_00253_),
    .Y(_00607_));
 sky130_fd_sc_hd__o211ai_4 _24895_ (.A1(_00242_),
    .A2(_00233_),
    .B1(_00253_),
    .C1(_00249_),
    .Y(_00608_));
 sky130_fd_sc_hd__o2111ai_4 _24896_ (.A1(net199),
    .A2(_00235_),
    .B1(_00603_),
    .C1(_00605_),
    .D1(_00608_),
    .Y(_00609_));
 sky130_fd_sc_hd__a22o_2 _24897_ (.A1(_00603_),
    .A2(_00605_),
    .B1(_00608_),
    .B2(_00239_),
    .X(_00610_));
 sky130_fd_sc_hd__o211ai_2 _24898_ (.A1(net270),
    .A2(net268),
    .B1(_00609_),
    .C1(_00610_),
    .Y(_00611_));
 sky130_fd_sc_hd__or3_1 _24899_ (.A(net270),
    .B(net268),
    .C(_00598_),
    .X(_00612_));
 sky130_fd_sc_hd__a21o_1 _24900_ (.A1(_00239_),
    .A2(_00608_),
    .B1(_00606_),
    .X(_00614_));
 sky130_fd_sc_hd__o21ai_1 _24901_ (.A1(_00243_),
    .A2(_00607_),
    .B1(_00606_),
    .Y(_00615_));
 sky130_fd_sc_hd__o311ai_2 _24902_ (.A1(_00243_),
    .A2(_00607_),
    .A3(_00606_),
    .B1(net244),
    .C1(_00615_),
    .Y(_00616_));
 sky130_fd_sc_hd__a31oi_4 _24903_ (.A1(_00610_),
    .A2(net244),
    .A3(_00609_),
    .B1(_00600_),
    .Y(_00617_));
 sky130_fd_sc_hd__a31o_4 _24904_ (.A1(_00610_),
    .A2(net244),
    .A3(_00609_),
    .B1(_00600_),
    .X(_00618_));
 sky130_fd_sc_hd__a311oi_1 _24905_ (.A1(_00610_),
    .A2(net244),
    .A3(_00609_),
    .B1(net200),
    .C1(_00600_),
    .Y(_00619_));
 sky130_fd_sc_hd__o211ai_4 _24906_ (.A1(net244),
    .A2(_00599_),
    .B1(_00611_),
    .C1(net198),
    .Y(_00620_));
 sky130_fd_sc_hd__a31oi_1 _24907_ (.A1(_00614_),
    .A2(_00615_),
    .A3(net244),
    .B1(net198),
    .Y(_00621_));
 sky130_fd_sc_hd__nand3_2 _24908_ (.A(_00616_),
    .B(net199),
    .C(_00612_),
    .Y(_00622_));
 sky130_fd_sc_hd__a21oi_2 _24909_ (.A1(_00621_),
    .A2(_00612_),
    .B1(_00619_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_2 _24910_ (.A(_00620_),
    .B(_00622_),
    .Y(_00625_));
 sky130_fd_sc_hd__and3_1 _24911_ (.A(_13510_),
    .B(_13947_),
    .C(_13948_),
    .X(_00626_));
 sky130_fd_sc_hd__o2111ai_4 _24912_ (.A1(_13507_),
    .A2(_13499_),
    .B1(_13505_),
    .C1(_13947_),
    .D1(_13948_),
    .Y(_00627_));
 sky130_fd_sc_hd__a211oi_4 _24913_ (.A1(_14325_),
    .A2(_14342_),
    .B1(_00627_),
    .C1(_14345_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand3_1 _24914_ (.A(_00268_),
    .B(_00626_),
    .C(_14347_),
    .Y(_00629_));
 sky130_fd_sc_hd__a32oi_2 _24915_ (.A1(_07936_),
    .A2(_00237_),
    .A3(_00260_),
    .B1(_00628_),
    .B2(_00268_),
    .Y(_00630_));
 sky130_fd_sc_hd__o211a_1 _24916_ (.A1(_00272_),
    .A2(_00267_),
    .B1(_00269_),
    .C1(_00629_),
    .X(_00631_));
 sky130_fd_sc_hd__o211ai_4 _24917_ (.A1(_00272_),
    .A2(_00267_),
    .B1(_00269_),
    .C1(_00629_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand3_2 _24918_ (.A(_00628_),
    .B(_00269_),
    .C(_00268_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand4_4 _24919_ (.A(_00628_),
    .B(_00269_),
    .C(_00268_),
    .D(_13521_),
    .Y(_00634_));
 sky130_fd_sc_hd__a2bb2oi_2 _24920_ (.A1_N(_13520_),
    .A2_N(_00633_),
    .B1(_00275_),
    .B2(_00630_),
    .Y(_00636_));
 sky130_fd_sc_hd__a21oi_1 _24921_ (.A1(_00632_),
    .A2(_00634_),
    .B1(_00625_),
    .Y(_00637_));
 sky130_fd_sc_hd__a21o_1 _24922_ (.A1(_00632_),
    .A2(_00634_),
    .B1(_00625_),
    .X(_00638_));
 sky130_fd_sc_hd__a31oi_2 _24923_ (.A1(_00625_),
    .A2(_00632_),
    .A3(_00634_),
    .B1(_05754_),
    .Y(_00639_));
 sky130_fd_sc_hd__a31o_1 _24924_ (.A1(_00625_),
    .A2(_00632_),
    .A3(_00634_),
    .B1(_05754_),
    .X(_00640_));
 sky130_fd_sc_hd__nand4_4 _24925_ (.A(_00620_),
    .B(_00622_),
    .C(_00632_),
    .D(_00634_),
    .Y(_00641_));
 sky130_fd_sc_hd__a22o_1 _24926_ (.A1(_00620_),
    .A2(_00622_),
    .B1(_00632_),
    .B2(_00634_),
    .X(_00642_));
 sky130_fd_sc_hd__o211a_1 _24927_ (.A1(net244),
    .A2(_00599_),
    .B1(_00611_),
    .C1(_05754_),
    .X(_00643_));
 sky130_fd_sc_hd__a311o_1 _24928_ (.A1(_00610_),
    .A2(net244),
    .A3(_00609_),
    .B1(net243),
    .C1(_00600_),
    .X(_00644_));
 sky130_fd_sc_hd__o221ai_4 _24929_ (.A1(net265),
    .A2(net264),
    .B1(_00623_),
    .B2(_00636_),
    .C1(_00641_),
    .Y(_00645_));
 sky130_fd_sc_hd__a22oi_4 _24930_ (.A1(_05754_),
    .A2(_00618_),
    .B1(_00639_),
    .B2(_00638_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2_2 _24931_ (.A(_05995_),
    .B(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__inv_2 _24932_ (.A(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__a311oi_4 _24933_ (.A1(_00642_),
    .A2(net243),
    .A3(_00641_),
    .B1(_00643_),
    .C1(_07936_),
    .Y(_00650_));
 sky130_fd_sc_hd__nand3_4 _24934_ (.A(_00645_),
    .B(_07935_),
    .C(_00644_),
    .Y(_00651_));
 sky130_fd_sc_hd__o221ai_4 _24935_ (.A1(net243),
    .A2(_00617_),
    .B1(_00637_),
    .B2(_00640_),
    .C1(_07936_),
    .Y(_00652_));
 sky130_fd_sc_hd__o221a_1 _24936_ (.A1(_14361_),
    .A2(_14366_),
    .B1(_00277_),
    .B2(_07564_),
    .C1(_14360_),
    .X(_00653_));
 sky130_fd_sc_hd__o211a_1 _24937_ (.A1(_14356_),
    .A2(net223),
    .B1(_00283_),
    .C1(_00279_),
    .X(_00654_));
 sky130_fd_sc_hd__a31o_1 _24938_ (.A1(_14362_),
    .A2(_00279_),
    .A3(_00283_),
    .B1(_00285_),
    .X(_00655_));
 sky130_fd_sc_hd__a31oi_4 _24939_ (.A1(_14362_),
    .A2(_00279_),
    .A3(_00283_),
    .B1(_00285_),
    .Y(_00656_));
 sky130_fd_sc_hd__a21oi_1 _24940_ (.A1(_00651_),
    .A2(_00652_),
    .B1(_00655_),
    .Y(_00658_));
 sky130_fd_sc_hd__o2bb2ai_4 _24941_ (.A1_N(_00651_),
    .A2_N(_00652_),
    .B1(_00653_),
    .B2(_00282_),
    .Y(_00659_));
 sky130_fd_sc_hd__o211a_1 _24942_ (.A1(_00285_),
    .A2(_00654_),
    .B1(_00652_),
    .C1(_00651_),
    .X(_00660_));
 sky130_fd_sc_hd__o211ai_4 _24943_ (.A1(_00285_),
    .A2(_00654_),
    .B1(_00652_),
    .C1(_00651_),
    .Y(_00661_));
 sky130_fd_sc_hd__a31oi_2 _24944_ (.A1(_00651_),
    .A2(_00652_),
    .A3(_00655_),
    .B1(_05995_),
    .Y(_00662_));
 sky130_fd_sc_hd__o211ai_4 _24945_ (.A1(net260),
    .A2(net255),
    .B1(_00659_),
    .C1(_00661_),
    .Y(_00663_));
 sky130_fd_sc_hd__o22ai_2 _24946_ (.A1(net260),
    .A2(net255),
    .B1(_00658_),
    .B2(_00660_),
    .Y(_00664_));
 sky130_fd_sc_hd__a31o_1 _24947_ (.A1(net240),
    .A2(_00659_),
    .A3(_00661_),
    .B1(_00649_),
    .X(_00665_));
 sky130_fd_sc_hd__o221ai_4 _24948_ (.A1(net227),
    .A2(_14375_),
    .B1(_07246_),
    .B2(_00294_),
    .C1(_14394_),
    .Y(_00666_));
 sky130_fd_sc_hd__o2bb2ai_1 _24949_ (.A1_N(_14377_),
    .A2_N(_14394_),
    .B1(_00293_),
    .B2(net223),
    .Y(_00667_));
 sky130_fd_sc_hd__a31o_1 _24950_ (.A1(net240),
    .A2(_00659_),
    .A3(_00661_),
    .B1(net202),
    .X(_00669_));
 sky130_fd_sc_hd__a211oi_4 _24951_ (.A1(_00662_),
    .A2(_00659_),
    .B1(_00649_),
    .C1(net202),
    .Y(_00670_));
 sky130_fd_sc_hd__nand3_2 _24952_ (.A(_00663_),
    .B(_07564_),
    .C(_00648_),
    .Y(_00671_));
 sky130_fd_sc_hd__a2bb2oi_4 _24953_ (.A1_N(net221),
    .A2_N(net220),
    .B1(_00648_),
    .B2(_00663_),
    .Y(_00672_));
 sky130_fd_sc_hd__o221ai_4 _24954_ (.A1(net221),
    .A2(net220),
    .B1(_00647_),
    .B2(net240),
    .C1(_00664_),
    .Y(_00673_));
 sky130_fd_sc_hd__nor2_1 _24955_ (.A(_00670_),
    .B(_00672_),
    .Y(_00674_));
 sky130_fd_sc_hd__o2111ai_1 _24956_ (.A1(_00294_),
    .A2(_07246_),
    .B1(_00671_),
    .C1(_00667_),
    .D1(_00673_),
    .Y(_00675_));
 sky130_fd_sc_hd__o2bb2ai_1 _24957_ (.A1_N(_00296_),
    .A2_N(_00667_),
    .B1(_00670_),
    .B2(_00672_),
    .Y(_00676_));
 sky130_fd_sc_hd__o2111ai_1 _24958_ (.A1(_00293_),
    .A2(net223),
    .B1(_00671_),
    .C1(_00666_),
    .D1(_00673_),
    .Y(_00677_));
 sky130_fd_sc_hd__o2bb2ai_1 _24959_ (.A1_N(_00297_),
    .A2_N(_00666_),
    .B1(_00670_),
    .B2(_00672_),
    .Y(_00678_));
 sky130_fd_sc_hd__nand3_2 _24960_ (.A(_00676_),
    .B(net214),
    .C(_00675_),
    .Y(_00680_));
 sky130_fd_sc_hd__a22o_1 _24961_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_00648_),
    .B2(_00663_),
    .X(_00681_));
 sky130_fd_sc_hd__nand3_2 _24962_ (.A(_00678_),
    .B(net214),
    .C(_00677_),
    .Y(_00682_));
 sky130_fd_sc_hd__o21a_1 _24963_ (.A1(net214),
    .A2(_00665_),
    .B1(_00680_),
    .X(_00683_));
 sky130_fd_sc_hd__o211ai_4 _24964_ (.A1(_07244_),
    .A2(net247),
    .B1(_00681_),
    .C1(_00682_),
    .Y(_00684_));
 sky130_fd_sc_hd__o211ai_4 _24965_ (.A1(_00665_),
    .A2(net214),
    .B1(net223),
    .C1(_00680_),
    .Y(_00685_));
 sky130_fd_sc_hd__nand2_1 _24966_ (.A(_00684_),
    .B(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__o2bb2ai_1 _24967_ (.A1_N(_00315_),
    .A2_N(_00316_),
    .B1(net227),
    .B2(_00308_),
    .Y(_00687_));
 sky130_fd_sc_hd__o211ai_2 _24968_ (.A1(net227),
    .A2(_00308_),
    .B1(_00320_),
    .C1(_00686_),
    .Y(_00688_));
 sky130_fd_sc_hd__o2111ai_4 _24969_ (.A1(_06924_),
    .A2(_00307_),
    .B1(_00684_),
    .C1(_00685_),
    .D1(_00687_),
    .Y(_00689_));
 sky130_fd_sc_hd__nand3_4 _24970_ (.A(_00689_),
    .B(net210),
    .C(_00688_),
    .Y(_00691_));
 sky130_fd_sc_hd__a211o_4 _24971_ (.A1(_00681_),
    .A2(_00682_),
    .B1(net238),
    .C1(_06610_),
    .X(_00692_));
 sky130_fd_sc_hd__nand2_2 _24972_ (.A(_00691_),
    .B(_00692_),
    .Y(_00693_));
 sky130_fd_sc_hd__inv_2 _24973_ (.A(_00693_),
    .Y(_00694_));
 sky130_fd_sc_hd__and3_1 _24974_ (.A(_06900_),
    .B(_06902_),
    .C(_00693_),
    .X(_00695_));
 sky130_fd_sc_hd__a211o_1 _24975_ (.A1(_00691_),
    .A2(_00692_),
    .B1(net231),
    .C1(net228),
    .X(_00696_));
 sky130_fd_sc_hd__a22oi_4 _24976_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_00691_),
    .B2(_00692_),
    .Y(_00697_));
 sky130_fd_sc_hd__a22o_2 _24977_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_00691_),
    .B2(_00692_),
    .X(_00698_));
 sky130_fd_sc_hd__and3_1 _24978_ (.A(_00691_),
    .B(_00692_),
    .C(_06922_),
    .X(_00699_));
 sky130_fd_sc_hd__o211ai_4 _24979_ (.A1(_06918_),
    .A2(_06920_),
    .B1(_00691_),
    .C1(_00692_),
    .Y(_00700_));
 sky130_fd_sc_hd__a41oi_2 _24980_ (.A1(_06915_),
    .A2(_06917_),
    .A3(_00691_),
    .A4(_00692_),
    .B1(_00697_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand4_2 _24981_ (.A(_13586_),
    .B(_13588_),
    .C(_14024_),
    .D(_14026_),
    .Y(_00703_));
 sky130_fd_sc_hd__a211oi_1 _24982_ (.A1(_14398_),
    .A2(_14416_),
    .B1(_00703_),
    .C1(_14419_),
    .Y(_00704_));
 sky130_fd_sc_hd__nand2_1 _24983_ (.A(_00331_),
    .B(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__o211ai_4 _24984_ (.A1(_00335_),
    .A2(_00330_),
    .B1(_00333_),
    .C1(_00705_),
    .Y(_00706_));
 sky130_fd_sc_hd__nor4b_2 _24985_ (.A(_14417_),
    .B(_00703_),
    .C(_14419_),
    .D_N(_13601_),
    .Y(_00707_));
 sky130_fd_sc_hd__o211ai_2 _24986_ (.A1(net235),
    .A2(_00325_),
    .B1(_00704_),
    .C1(_13601_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand3_4 _24987_ (.A(_00331_),
    .B(_00333_),
    .C(_00707_),
    .Y(_00709_));
 sky130_fd_sc_hd__o21ai_4 _24988_ (.A1(_00330_),
    .A2(_00708_),
    .B1(_00706_),
    .Y(_00710_));
 sky130_fd_sc_hd__o211ai_1 _24989_ (.A1(_00697_),
    .A2(_00699_),
    .B1(_00706_),
    .C1(_00709_),
    .Y(_00711_));
 sky130_fd_sc_hd__nand2_1 _24990_ (.A(_00710_),
    .B(_00702_),
    .Y(_00713_));
 sky130_fd_sc_hd__a22o_1 _24991_ (.A1(_00698_),
    .A2(_00700_),
    .B1(_00706_),
    .B2(_00709_),
    .X(_00714_));
 sky130_fd_sc_hd__o211ai_1 _24992_ (.A1(_06924_),
    .A2(_00693_),
    .B1(_00706_),
    .C1(_00709_),
    .Y(_00715_));
 sky130_fd_sc_hd__nand4_4 _24993_ (.A(_00698_),
    .B(_00700_),
    .C(_00706_),
    .D(_00709_),
    .Y(_00716_));
 sky130_fd_sc_hd__nand3_1 _24994_ (.A(_00714_),
    .B(_00716_),
    .C(net208),
    .Y(_00717_));
 sky130_fd_sc_hd__nand3_1 _24995_ (.A(_00713_),
    .B(net208),
    .C(_00711_),
    .Y(_00718_));
 sky130_fd_sc_hd__o211a_2 _24996_ (.A1(net208),
    .A2(_00693_),
    .B1(_07232_),
    .C1(_00718_),
    .X(_00719_));
 sky130_fd_sc_hd__a211o_1 _24997_ (.A1(_00696_),
    .A2(_00717_),
    .B1(net207),
    .C1(net205),
    .X(_00720_));
 sky130_fd_sc_hd__a31o_1 _24998_ (.A1(_00714_),
    .A2(_00716_),
    .A3(net208),
    .B1(net233),
    .X(_00721_));
 sky130_fd_sc_hd__a311oi_2 _24999_ (.A1(_00714_),
    .A2(_00716_),
    .A3(net208),
    .B1(_00695_),
    .C1(net233),
    .Y(_00722_));
 sky130_fd_sc_hd__nand3_4 _25000_ (.A(_00717_),
    .B(net235),
    .C(_00696_),
    .Y(_00724_));
 sky130_fd_sc_hd__o211ai_4 _25001_ (.A1(_00693_),
    .A2(net208),
    .B1(net233),
    .C1(_00718_),
    .Y(_00725_));
 sky130_fd_sc_hd__a21oi_1 _25002_ (.A1(net252),
    .A2(_00343_),
    .B1(_00346_),
    .Y(_00726_));
 sky130_fd_sc_hd__o32a_2 _25003_ (.A1(net284),
    .A2(net282),
    .A3(_00343_),
    .B1(_00346_),
    .B2(_00351_),
    .X(_00727_));
 sky130_fd_sc_hd__a21oi_1 _25004_ (.A1(_00349_),
    .A2(_00346_),
    .B1(_00351_),
    .Y(_00728_));
 sky130_fd_sc_hd__a21oi_1 _25005_ (.A1(_00724_),
    .A2(_00725_),
    .B1(_00727_),
    .Y(_00729_));
 sky130_fd_sc_hd__o2bb2ai_4 _25006_ (.A1_N(_00724_),
    .A2_N(_00725_),
    .B1(_00726_),
    .B2(_00348_),
    .Y(_00730_));
 sky130_fd_sc_hd__o211a_1 _25007_ (.A1(_00695_),
    .A2(_00721_),
    .B1(_00725_),
    .C1(_00727_),
    .X(_00731_));
 sky130_fd_sc_hd__o211ai_2 _25008_ (.A1(_00695_),
    .A2(_00721_),
    .B1(_00725_),
    .C1(_00727_),
    .Y(_00732_));
 sky130_fd_sc_hd__a31oi_4 _25009_ (.A1(_00727_),
    .A2(_00725_),
    .A3(_00724_),
    .B1(_07232_),
    .Y(_00733_));
 sky130_fd_sc_hd__o211ai_2 _25010_ (.A1(net207),
    .A2(net205),
    .B1(_00730_),
    .C1(_00732_),
    .Y(_00735_));
 sky130_fd_sc_hd__a311o_1 _25011_ (.A1(_00714_),
    .A2(_00716_),
    .A3(net208),
    .B1(_07233_),
    .C1(_00695_),
    .X(_00736_));
 sky130_fd_sc_hd__o22ai_2 _25012_ (.A1(net207),
    .A2(net205),
    .B1(_00729_),
    .B2(_00731_),
    .Y(_00737_));
 sky130_fd_sc_hd__a31o_1 _25013_ (.A1(_07233_),
    .A2(_00730_),
    .A3(_00732_),
    .B1(_00719_),
    .X(_00738_));
 sky130_fd_sc_hd__o311a_1 _25014_ (.A1(_05765_),
    .A2(net288),
    .A3(_14448_),
    .B1(_00003_),
    .C1(_00364_),
    .X(_00739_));
 sky130_fd_sc_hd__o2bb2ai_1 _25015_ (.A1_N(_14450_),
    .A2_N(_00003_),
    .B1(_00362_),
    .B2(_06014_),
    .Y(_00740_));
 sky130_fd_sc_hd__o32a_1 _25016_ (.A1(_06009_),
    .A2(net287),
    .A3(_00362_),
    .B1(_00363_),
    .B2(_00369_),
    .X(_00741_));
 sky130_fd_sc_hd__o32ai_4 _25017_ (.A1(_06009_),
    .A2(net287),
    .A3(_00362_),
    .B1(_00363_),
    .B2(_00369_),
    .Y(_00742_));
 sky130_fd_sc_hd__a21oi_1 _25018_ (.A1(_00733_),
    .A2(_00730_),
    .B1(net252),
    .Y(_00743_));
 sky130_fd_sc_hd__o2bb2ai_1 _25019_ (.A1_N(_00730_),
    .A2_N(_00733_),
    .B1(_06309_),
    .B2(_06312_),
    .Y(_00744_));
 sky130_fd_sc_hd__a211oi_4 _25020_ (.A1(_00733_),
    .A2(_00730_),
    .B1(_00719_),
    .C1(net252),
    .Y(_00746_));
 sky130_fd_sc_hd__a2bb2oi_2 _25021_ (.A1_N(net284),
    .A2_N(net282),
    .B1(_00720_),
    .B2(_00735_),
    .Y(_00747_));
 sky130_fd_sc_hd__o211ai_4 _25022_ (.A1(net284),
    .A2(net282),
    .B1(_00736_),
    .C1(_00737_),
    .Y(_00748_));
 sky130_fd_sc_hd__o211ai_1 _25023_ (.A1(_00744_),
    .A2(_00719_),
    .B1(_00742_),
    .C1(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__o2bb2ai_1 _25024_ (.A1_N(_00364_),
    .A2_N(_00740_),
    .B1(_00746_),
    .B2(_00747_),
    .Y(_00750_));
 sky130_fd_sc_hd__nand3_2 _25025_ (.A(_00750_),
    .B(net163),
    .C(_00749_),
    .Y(_00751_));
 sky130_fd_sc_hd__and3_1 _25026_ (.A(_07550_),
    .B(_00736_),
    .C(_00737_),
    .X(_00752_));
 sky130_fd_sc_hd__a211o_1 _25027_ (.A1(_00720_),
    .A2(_00735_),
    .B1(_07544_),
    .C1(_07546_),
    .X(_00753_));
 sky130_fd_sc_hd__o211ai_2 _25028_ (.A1(_00719_),
    .A2(_00744_),
    .B1(_00748_),
    .C1(_00741_),
    .Y(_00754_));
 sky130_fd_sc_hd__o22ai_2 _25029_ (.A1(_00365_),
    .A2(_00739_),
    .B1(_00746_),
    .B2(_00747_),
    .Y(_00755_));
 sky130_fd_sc_hd__nand3_1 _25030_ (.A(_00754_),
    .B(_00755_),
    .C(net163),
    .Y(_00757_));
 sky130_fd_sc_hd__a31oi_2 _25031_ (.A1(_00754_),
    .A2(_00755_),
    .A3(net163),
    .B1(_00752_),
    .Y(_00758_));
 sky130_fd_sc_hd__o211a_1 _25032_ (.A1(_00738_),
    .A2(net163),
    .B1(_06014_),
    .C1(_00751_),
    .X(_00759_));
 sky130_fd_sc_hd__o211ai_4 _25033_ (.A1(_00738_),
    .A2(net163),
    .B1(_06014_),
    .C1(_00751_),
    .Y(_00760_));
 sky130_fd_sc_hd__and3_1 _25034_ (.A(_00757_),
    .B(net254),
    .C(_00753_),
    .X(_00761_));
 sky130_fd_sc_hd__nand3_4 _25035_ (.A(_00757_),
    .B(net254),
    .C(_00753_),
    .Y(_00762_));
 sky130_fd_sc_hd__a2bb2oi_1 _25036_ (.A1_N(net263),
    .A2_N(_00376_),
    .B1(_00384_),
    .B2(_00012_),
    .Y(_00763_));
 sky130_fd_sc_hd__o21ai_2 _25037_ (.A1(net263),
    .A2(_00376_),
    .B1(_00386_),
    .Y(_00764_));
 sky130_fd_sc_hd__o2bb2ai_4 _25038_ (.A1_N(_00760_),
    .A2_N(_00762_),
    .B1(_00763_),
    .B2(_00381_),
    .Y(_00765_));
 sky130_fd_sc_hd__nand4_4 _25039_ (.A(_00382_),
    .B(_00760_),
    .C(_00762_),
    .D(_00764_),
    .Y(_00766_));
 sky130_fd_sc_hd__nand3_4 _25040_ (.A(_00765_),
    .B(_00766_),
    .C(net162),
    .Y(_00768_));
 sky130_fd_sc_hd__o211a_1 _25041_ (.A1(_00738_),
    .A2(net163),
    .B1(_07917_),
    .C1(_00751_),
    .X(_00769_));
 sky130_fd_sc_hd__or3_4 _25042_ (.A(net183),
    .B(net182),
    .C(_00758_),
    .X(_00770_));
 sky130_fd_sc_hd__a31oi_2 _25043_ (.A1(_00765_),
    .A2(_00766_),
    .A3(net162),
    .B1(_00769_),
    .Y(_00771_));
 sky130_fd_sc_hd__a21oi_4 _25044_ (.A1(_00768_),
    .A2(_00770_),
    .B1(net159),
    .Y(_00772_));
 sky130_fd_sc_hd__inv_2 _25045_ (.A(_00772_),
    .Y(_00773_));
 sky130_fd_sc_hd__a21oi_4 _25046_ (.A1(_00768_),
    .A2(_00770_),
    .B1(net263),
    .Y(_00774_));
 sky130_fd_sc_hd__a22o_2 _25047_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_00768_),
    .B2(_00770_),
    .X(_00775_));
 sky130_fd_sc_hd__a31oi_1 _25048_ (.A1(_00765_),
    .A2(_00766_),
    .A3(net162),
    .B1(_05768_),
    .Y(_00776_));
 sky130_fd_sc_hd__o221a_1 _25049_ (.A1(_05765_),
    .A2(net288),
    .B1(net161),
    .B2(_00758_),
    .C1(_00768_),
    .X(_00777_));
 sky130_fd_sc_hd__a311o_2 _25050_ (.A1(_00765_),
    .A2(_00766_),
    .A3(net162),
    .B1(_00769_),
    .C1(_05768_),
    .X(_00779_));
 sky130_fd_sc_hd__a21oi_1 _25051_ (.A1(_00770_),
    .A2(_00776_),
    .B1(_00774_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand4_2 _25052_ (.A(_13665_),
    .B(_13667_),
    .C(_14097_),
    .D(_14099_),
    .Y(_00781_));
 sky130_fd_sc_hd__a21oi_2 _25053_ (.A1(net294),
    .A2(_00026_),
    .B1(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__nor3_1 _25054_ (.A(_00032_),
    .B(_00781_),
    .C(_00035_),
    .Y(_00783_));
 sky130_fd_sc_hd__o211ai_2 _25055_ (.A1(net294),
    .A2(_00026_),
    .B1(_00782_),
    .C1(_00399_),
    .Y(_00784_));
 sky130_fd_sc_hd__o211a_1 _25056_ (.A1(_00404_),
    .A2(_00398_),
    .B1(_00400_),
    .C1(_00784_),
    .X(_00785_));
 sky130_fd_sc_hd__o211ai_4 _25057_ (.A1(_00404_),
    .A2(_00398_),
    .B1(_00400_),
    .C1(_00784_),
    .Y(_00786_));
 sky130_fd_sc_hd__o211ai_1 _25058_ (.A1(net294),
    .A2(_00026_),
    .B1(_00782_),
    .C1(_13678_),
    .Y(_00787_));
 sky130_fd_sc_hd__nand4_4 _25059_ (.A(_00782_),
    .B(_00400_),
    .C(_00399_),
    .D(_00034_),
    .Y(_00788_));
 sky130_fd_sc_hd__nand4_1 _25060_ (.A(_00399_),
    .B(_00783_),
    .C(_00400_),
    .D(_13678_),
    .Y(_00790_));
 sky130_fd_sc_hd__o21ai_1 _25061_ (.A1(_13680_),
    .A2(_00788_),
    .B1(_00786_),
    .Y(_00791_));
 sky130_fd_sc_hd__and3_1 _25062_ (.A(_00775_),
    .B(_00779_),
    .C(_00791_),
    .X(_00792_));
 sky130_fd_sc_hd__nand2_1 _25063_ (.A(_00791_),
    .B(_00780_),
    .Y(_00793_));
 sky130_fd_sc_hd__o221ai_2 _25064_ (.A1(_13680_),
    .A2(_00788_),
    .B1(_00777_),
    .B2(_00774_),
    .C1(_00786_),
    .Y(_00794_));
 sky130_fd_sc_hd__a22o_2 _25065_ (.A1(_00775_),
    .A2(_00779_),
    .B1(_00786_),
    .B2(_00790_),
    .X(_00795_));
 sky130_fd_sc_hd__o2bb2ai_1 _25066_ (.A1_N(net263),
    .A2_N(_00771_),
    .B1(_00787_),
    .B2(_00401_),
    .Y(_00796_));
 sky130_fd_sc_hd__o211ai_4 _25067_ (.A1(_13680_),
    .A2(_00788_),
    .B1(_00786_),
    .C1(_00779_),
    .Y(_00797_));
 sky130_fd_sc_hd__o2111ai_4 _25068_ (.A1(_13680_),
    .A2(_00788_),
    .B1(_00786_),
    .C1(_00779_),
    .D1(_00775_),
    .Y(_00798_));
 sky130_fd_sc_hd__a22oi_2 _25069_ (.A1(_08297_),
    .A2(_08299_),
    .B1(_00793_),
    .B2(_00794_),
    .Y(_00799_));
 sky130_fd_sc_hd__o221ai_4 _25070_ (.A1(_08296_),
    .A2(net179),
    .B1(_00774_),
    .B2(_00797_),
    .C1(_00795_),
    .Y(_00801_));
 sky130_fd_sc_hd__a31oi_4 _25071_ (.A1(_00795_),
    .A2(_00798_),
    .A3(net159),
    .B1(_00772_),
    .Y(_00802_));
 sky130_fd_sc_hd__o22a_2 _25072_ (.A1(_08705_),
    .A2(_08707_),
    .B1(_00772_),
    .B2(_00799_),
    .X(_00803_));
 sky130_fd_sc_hd__or3_1 _25073_ (.A(net158),
    .B(_08712_),
    .C(_00802_),
    .X(_00804_));
 sky130_fd_sc_hd__a31o_2 _25074_ (.A1(_00795_),
    .A2(_00798_),
    .A3(net159),
    .B1(net292),
    .X(_00805_));
 sky130_fd_sc_hd__a311oi_4 _25075_ (.A1(_00795_),
    .A2(_00798_),
    .A3(net159),
    .B1(_00772_),
    .C1(net292),
    .Y(_00806_));
 sky130_fd_sc_hd__a311o_2 _25076_ (.A1(_00795_),
    .A2(_00798_),
    .A3(net159),
    .B1(_00772_),
    .C1(net292),
    .X(_00807_));
 sky130_fd_sc_hd__a2bb2oi_4 _25077_ (.A1_N(_05500_),
    .A2_N(_05503_),
    .B1(_00773_),
    .B2(_00801_),
    .Y(_00808_));
 sky130_fd_sc_hd__o22ai_2 _25078_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_00772_),
    .B2(_00799_),
    .Y(_00809_));
 sky130_fd_sc_hd__o32a_4 _25079_ (.A1(net318),
    .A2(net315),
    .A3(_00410_),
    .B1(_00413_),
    .B2(_00417_),
    .X(_00810_));
 sky130_fd_sc_hd__o31a_1 _25080_ (.A1(_00048_),
    .A2(_00411_),
    .A3(_00415_),
    .B1(_00418_),
    .X(_00812_));
 sky130_fd_sc_hd__o21a_1 _25081_ (.A1(_00806_),
    .A2(_00808_),
    .B1(_00812_),
    .X(_00813_));
 sky130_fd_sc_hd__o21ai_4 _25082_ (.A1(_00806_),
    .A2(_00808_),
    .B1(_00812_),
    .Y(_00814_));
 sky130_fd_sc_hd__o21ai_1 _25083_ (.A1(_05507_),
    .A2(_00802_),
    .B1(_00810_),
    .Y(_00815_));
 sky130_fd_sc_hd__o211ai_4 _25084_ (.A1(_00772_),
    .A2(_00805_),
    .B1(_00810_),
    .C1(_00809_),
    .Y(_00816_));
 sky130_fd_sc_hd__o22ai_2 _25085_ (.A1(_08709_),
    .A2(_08712_),
    .B1(_00806_),
    .B2(_00815_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand3_2 _25086_ (.A(_00814_),
    .B(_00816_),
    .C(net149),
    .Y(_00818_));
 sky130_fd_sc_hd__a31oi_4 _25087_ (.A1(_00814_),
    .A2(_00816_),
    .A3(net149),
    .B1(_00803_),
    .Y(_00819_));
 sky130_fd_sc_hd__o22ai_4 _25088_ (.A1(net149),
    .A2(_00802_),
    .B1(_00813_),
    .B2(_00817_),
    .Y(_00820_));
 sky130_fd_sc_hd__a311o_1 _25089_ (.A1(_00814_),
    .A2(_00816_),
    .A3(net149),
    .B1(net146),
    .C1(_00803_),
    .X(_00821_));
 sky130_fd_sc_hd__and3_1 _25090_ (.A(_00062_),
    .B(_00075_),
    .C(_00429_),
    .X(_00823_));
 sky130_fd_sc_hd__a31oi_2 _25091_ (.A1(_00062_),
    .A2(_00075_),
    .A3(_00429_),
    .B1(_00430_),
    .Y(_00824_));
 sky130_fd_sc_hd__a31o_1 _25092_ (.A1(_00062_),
    .A2(_00075_),
    .A3(_00429_),
    .B1(_00430_),
    .X(_00825_));
 sky130_fd_sc_hd__a311oi_2 _25093_ (.A1(_00814_),
    .A2(_00816_),
    .A3(net149),
    .B1(_00803_),
    .C1(_05249_),
    .Y(_00826_));
 sky130_fd_sc_hd__o211ai_4 _25094_ (.A1(net149),
    .A2(_00802_),
    .B1(_05248_),
    .C1(_00818_),
    .Y(_00827_));
 sky130_fd_sc_hd__a2bb2oi_1 _25095_ (.A1_N(net318),
    .A2_N(net315),
    .B1(_00804_),
    .B2(_00818_),
    .Y(_00828_));
 sky130_fd_sc_hd__o21ai_2 _25096_ (.A1(net318),
    .A2(net315),
    .B1(_00820_),
    .Y(_00829_));
 sky130_fd_sc_hd__o211ai_1 _25097_ (.A1(_00430_),
    .A2(_00823_),
    .B1(_00827_),
    .C1(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__o21ai_1 _25098_ (.A1(_00826_),
    .A2(_00828_),
    .B1(_00824_),
    .Y(_00831_));
 sky130_fd_sc_hd__o211ai_2 _25099_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_00830_),
    .C1(_00831_),
    .Y(_00832_));
 sky130_fd_sc_hd__a21oi_2 _25100_ (.A1(_00804_),
    .A2(_00818_),
    .B1(net146),
    .Y(_00834_));
 sky130_fd_sc_hd__nand3_1 _25101_ (.A(_00829_),
    .B(_00824_),
    .C(_00827_),
    .Y(_00835_));
 sky130_fd_sc_hd__o22ai_2 _25102_ (.A1(_00430_),
    .A2(_00823_),
    .B1(_00826_),
    .B2(_00828_),
    .Y(_00836_));
 sky130_fd_sc_hd__o211ai_2 _25103_ (.A1(_09120_),
    .A2(_09121_),
    .B1(_00835_),
    .C1(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hd__a31o_1 _25104_ (.A1(net146),
    .A2(_00835_),
    .A3(_00836_),
    .B1(_00834_),
    .X(_00838_));
 sky130_fd_sc_hd__o31a_2 _25105_ (.A1(_09120_),
    .A2(_09121_),
    .A3(_00819_),
    .B1(_00837_),
    .X(_00839_));
 sky130_fd_sc_hd__o211ai_4 _25106_ (.A1(net340),
    .A2(_04184_),
    .B1(_00821_),
    .C1(_00832_),
    .Y(_00840_));
 sky130_fd_sc_hd__a31o_1 _25107_ (.A1(net146),
    .A2(_00835_),
    .A3(_00836_),
    .B1(_04238_),
    .X(_00841_));
 sky130_fd_sc_hd__o211ai_4 _25108_ (.A1(net146),
    .A2(_00819_),
    .B1(_04227_),
    .C1(_00837_),
    .Y(_00842_));
 sky130_fd_sc_hd__a31o_1 _25109_ (.A1(_00447_),
    .A2(_00455_),
    .A3(_00457_),
    .B1(_00444_),
    .X(_00843_));
 sky130_fd_sc_hd__a31oi_2 _25110_ (.A1(_00447_),
    .A2(_00455_),
    .A3(_00457_),
    .B1(_00444_),
    .Y(_00845_));
 sky130_fd_sc_hd__o2111ai_1 _25111_ (.A1(_02137_),
    .A2(_00442_),
    .B1(_00461_),
    .C1(_00840_),
    .D1(_00842_),
    .Y(_00846_));
 sky130_fd_sc_hd__a22o_1 _25112_ (.A1(_00445_),
    .A2(_00461_),
    .B1(_00840_),
    .B2(_00842_),
    .X(_00847_));
 sky130_fd_sc_hd__o211ai_2 _25113_ (.A1(_09553_),
    .A2(net155),
    .B1(_00846_),
    .C1(_00847_),
    .Y(_00848_));
 sky130_fd_sc_hd__a21oi_2 _25114_ (.A1(_00840_),
    .A2(_00842_),
    .B1(_00843_),
    .Y(_00849_));
 sky130_fd_sc_hd__a31o_1 _25115_ (.A1(_00843_),
    .A2(_00842_),
    .A3(_00840_),
    .B1(_09562_),
    .X(_00850_));
 sky130_fd_sc_hd__o22ai_4 _25116_ (.A1(net143),
    .A2(_00839_),
    .B1(_00849_),
    .B2(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__o211a_2 _25117_ (.A1(_00838_),
    .A2(net143),
    .B1(_02148_),
    .C1(_00848_),
    .X(_00852_));
 sky130_fd_sc_hd__o2111ai_4 _25118_ (.A1(_00838_),
    .A2(net143),
    .B1(_02126_),
    .C1(_02104_),
    .D1(_00848_),
    .Y(_00853_));
 sky130_fd_sc_hd__o221ai_4 _25119_ (.A1(net143),
    .A2(_00839_),
    .B1(_00849_),
    .B2(_00850_),
    .C1(_02137_),
    .Y(_00854_));
 sky130_fd_sc_hd__o2111ai_2 _25120_ (.A1(_13742_),
    .A2(_13736_),
    .B1(_13741_),
    .C1(_14161_),
    .D1(_14164_),
    .Y(_00856_));
 sky130_fd_sc_hd__a21oi_1 _25121_ (.A1(_12899_),
    .A2(_00095_),
    .B1(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__nor3_1 _25122_ (.A(_00856_),
    .B(_00101_),
    .C(_00099_),
    .Y(_00858_));
 sky130_fd_sc_hd__o211ai_2 _25123_ (.A1(_12899_),
    .A2(_00095_),
    .B1(_00857_),
    .C1(_00472_),
    .Y(_00859_));
 sky130_fd_sc_hd__o211ai_4 _25124_ (.A1(_00477_),
    .A2(_00470_),
    .B1(_00474_),
    .C1(_00859_),
    .Y(_00860_));
 sky130_fd_sc_hd__nand4_4 _25125_ (.A(_00472_),
    .B(_00858_),
    .C(_00474_),
    .D(_13744_),
    .Y(_00861_));
 sky130_fd_sc_hd__nand2_1 _25126_ (.A(_00860_),
    .B(_00861_),
    .Y(_00862_));
 sky130_fd_sc_hd__a22oi_1 _25127_ (.A1(_00853_),
    .A2(_00854_),
    .B1(_00860_),
    .B2(_00861_),
    .Y(_00863_));
 sky130_fd_sc_hd__a22o_1 _25128_ (.A1(_00853_),
    .A2(_00854_),
    .B1(_00860_),
    .B2(_00861_),
    .X(_00864_));
 sky130_fd_sc_hd__o211ai_2 _25129_ (.A1(_00851_),
    .A2(_02148_),
    .B1(_00861_),
    .C1(_00860_),
    .Y(_00865_));
 sky130_fd_sc_hd__o2111a_1 _25130_ (.A1(_02148_),
    .A2(_00851_),
    .B1(_00853_),
    .C1(_00860_),
    .D1(_00861_),
    .X(_00867_));
 sky130_fd_sc_hd__o221ai_4 _25131_ (.A1(_09571_),
    .A2(_09573_),
    .B1(_00852_),
    .B2(_00865_),
    .C1(_00864_),
    .Y(_00868_));
 sky130_fd_sc_hd__nand2_1 _25132_ (.A(_09578_),
    .B(_00851_),
    .Y(_00869_));
 sky130_fd_sc_hd__a211o_2 _25133_ (.A1(_00868_),
    .A2(_00869_),
    .B1(_10474_),
    .C1(net138),
    .X(_00870_));
 sky130_fd_sc_hd__inv_2 _25134_ (.A(_00870_),
    .Y(_00871_));
 sky130_fd_sc_hd__o311a_1 _25135_ (.A1(_09578_),
    .A2(_00863_),
    .A3(_00867_),
    .B1(_00869_),
    .C1(_00240_),
    .X(_00872_));
 sky130_fd_sc_hd__nand3_2 _25136_ (.A(_00868_),
    .B(_00869_),
    .C(_00240_),
    .Y(_00873_));
 sky130_fd_sc_hd__a21oi_1 _25137_ (.A1(_00868_),
    .A2(_00869_),
    .B1(_00240_),
    .Y(_00874_));
 sky130_fd_sc_hd__a22o_2 _25138_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_00868_),
    .B2(_00869_),
    .X(_00875_));
 sky130_fd_sc_hd__a21oi_2 _25139_ (.A1(_00484_),
    .A2(_00486_),
    .B1(_00487_),
    .Y(_00876_));
 sky130_fd_sc_hd__o21ai_1 _25140_ (.A1(_00872_),
    .A2(_00874_),
    .B1(_00876_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand3b_1 _25141_ (.A_N(_00876_),
    .B(_00875_),
    .C(_00873_),
    .Y(_00879_));
 sky130_fd_sc_hd__o311a_1 _25142_ (.A1(_00872_),
    .A2(_00876_),
    .A3(_00874_),
    .B1(net131),
    .C1(_00878_),
    .X(_00880_));
 sky130_fd_sc_hd__nand3_1 _25143_ (.A(net131),
    .B(_00878_),
    .C(_00879_),
    .Y(_00881_));
 sky130_fd_sc_hd__nor2_1 _25144_ (.A(_00871_),
    .B(_00880_),
    .Y(_00882_));
 sky130_fd_sc_hd__a31oi_1 _25145_ (.A1(net131),
    .A2(_00878_),
    .A3(_00879_),
    .B1(_12899_),
    .Y(_00883_));
 sky130_fd_sc_hd__o211a_1 _25146_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_00870_),
    .C1(_00881_),
    .X(_00884_));
 sky130_fd_sc_hd__a2bb2oi_1 _25147_ (.A1_N(net361),
    .A2_N(net345),
    .B1(_00870_),
    .B2(_00881_),
    .Y(_00885_));
 sky130_fd_sc_hd__o21ai_1 _25148_ (.A1(_00871_),
    .A2(_00880_),
    .B1(_12899_),
    .Y(_00886_));
 sky130_fd_sc_hd__a21oi_1 _25149_ (.A1(_00870_),
    .A2(_00883_),
    .B1(_00885_),
    .Y(_00887_));
 sky130_fd_sc_hd__a21oi_1 _25150_ (.A1(_00494_),
    .A2(_00496_),
    .B1(_00497_),
    .Y(_00889_));
 sky130_fd_sc_hd__o21ai_1 _25151_ (.A1(_00884_),
    .A2(_00885_),
    .B1(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__a31oi_2 _25152_ (.A1(_00870_),
    .A2(_00881_),
    .A3(_12888_),
    .B1(_00889_),
    .Y(_00891_));
 sky130_fd_sc_hd__a21oi_1 _25153_ (.A1(_00891_),
    .A2(_00886_),
    .B1(_10953_),
    .Y(_00892_));
 sky130_fd_sc_hd__o2bb2ai_2 _25154_ (.A1_N(_00890_),
    .A2_N(_00892_),
    .B1(_10954_),
    .B2(_00882_),
    .Y(_00893_));
 sky130_fd_sc_hd__o2bb2a_1 _25155_ (.A1_N(_00890_),
    .A2_N(_00892_),
    .B1(_10954_),
    .B2(_00882_),
    .X(_00894_));
 sky130_fd_sc_hd__a21oi_2 _25156_ (.A1(_00506_),
    .A2(_00508_),
    .B1(_00505_),
    .Y(_00895_));
 sky130_fd_sc_hd__a21oi_2 _25157_ (.A1(_11265_),
    .A2(_11287_),
    .B1(_00893_),
    .Y(_00896_));
 sky130_fd_sc_hd__and3_1 _25158_ (.A(_00893_),
    .B(_11287_),
    .C(_11265_),
    .X(_00897_));
 sky130_fd_sc_hd__o21ai_1 _25159_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_00893_),
    .Y(_00898_));
 sky130_fd_sc_hd__a31o_1 _25160_ (.A1(_11265_),
    .A2(_11287_),
    .A3(_00893_),
    .B1(_00895_),
    .X(_00900_));
 sky130_fd_sc_hd__o21ai_1 _25161_ (.A1(_00896_),
    .A2(_00897_),
    .B1(_00895_),
    .Y(_00901_));
 sky130_fd_sc_hd__o211ai_2 _25162_ (.A1(_00896_),
    .A2(_00900_),
    .B1(_00901_),
    .C1(_11465_),
    .Y(_00902_));
 sky130_fd_sc_hd__o21ai_2 _25163_ (.A1(_11465_),
    .A2(_00894_),
    .B1(_00902_),
    .Y(_00903_));
 sky130_fd_sc_hd__and3_1 _25164_ (.A(_00903_),
    .B(_10004_),
    .C(_09982_),
    .X(_00904_));
 sky130_fd_sc_hd__o221a_1 _25165_ (.A1(net365),
    .A2(net362),
    .B1(_11465_),
    .B2(_00894_),
    .C1(_00902_),
    .X(_00905_));
 sky130_fd_sc_hd__a32o_1 _25166_ (.A1(_08918_),
    .A2(_00503_),
    .A3(_00510_),
    .B1(_00513_),
    .B2(_00516_),
    .X(_00906_));
 sky130_fd_sc_hd__o21bai_1 _25167_ (.A1(_00904_),
    .A2(_00905_),
    .B1_N(_00906_),
    .Y(_00907_));
 sky130_fd_sc_hd__a21o_1 _25168_ (.A1(_00907_),
    .A2(_11943_),
    .B1(_00903_),
    .X(_00908_));
 sky130_fd_sc_hd__and3_1 _25169_ (.A(_05119_),
    .B(_00521_),
    .C(_00908_),
    .X(_00909_));
 sky130_fd_sc_hd__a21oi_1 _25170_ (.A1(_05119_),
    .A2(_00521_),
    .B1(_00908_),
    .Y(_00911_));
 sky130_fd_sc_hd__nor2_1 _25171_ (.A(_00909_),
    .B(_00911_),
    .Y(net97));
 sky130_fd_sc_hd__o21ai_1 _25172_ (.A1(_00908_),
    .A2(_00521_),
    .B1(_05119_),
    .Y(_00912_));
 sky130_fd_sc_hd__o211ai_1 _25173_ (.A1(_00523_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_00532_),
    .Y(_00913_));
 sky130_fd_sc_hd__a311o_2 _25174_ (.A1(_11471_),
    .A2(_00526_),
    .A3(_00532_),
    .B1(net308),
    .C1(_12703_),
    .X(_00914_));
 sky130_fd_sc_hd__and3_1 _25175_ (.A(_00913_),
    .B(net311),
    .C(_10971_),
    .X(_00915_));
 sky130_fd_sc_hd__a311o_1 _25176_ (.A1(_11471_),
    .A2(_00526_),
    .A3(_00532_),
    .B1(_10970_),
    .C1(_12703_),
    .X(_00916_));
 sky130_fd_sc_hd__o2bb2a_1 _25177_ (.A1_N(net311),
    .A2_N(_00913_),
    .B1(_10967_),
    .B2(_10965_),
    .X(_00917_));
 sky130_fd_sc_hd__nor2_1 _25178_ (.A(_00915_),
    .B(_00917_),
    .Y(_00918_));
 sky130_fd_sc_hd__o21ai_1 _25179_ (.A1(_00541_),
    .A2(_00544_),
    .B1(_00540_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand2_1 _25180_ (.A(_00919_),
    .B(_00918_),
    .Y(_00921_));
 sky130_fd_sc_hd__o221ai_4 _25181_ (.A1(_00541_),
    .A2(_00544_),
    .B1(_00915_),
    .B2(_00917_),
    .C1(_00540_),
    .Y(_00922_));
 sky130_fd_sc_hd__nand3_2 _25182_ (.A(_00921_),
    .B(_00922_),
    .C(net307),
    .Y(_00923_));
 sky130_fd_sc_hd__and2_1 _25183_ (.A(_00914_),
    .B(_00923_),
    .X(_00924_));
 sky130_fd_sc_hd__a21oi_4 _25184_ (.A1(_00914_),
    .A2(_00923_),
    .B1(net278),
    .Y(_00925_));
 sky130_fd_sc_hd__a2bb2oi_1 _25185_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_00914_),
    .B2(_00923_),
    .Y(_00926_));
 sky130_fd_sc_hd__a31oi_1 _25186_ (.A1(_00921_),
    .A2(_00922_),
    .A3(net307),
    .B1(_10492_),
    .Y(_00927_));
 sky130_fd_sc_hd__and3_1 _25187_ (.A(_00923_),
    .B(net150),
    .C(_00914_),
    .X(_00928_));
 sky130_fd_sc_hd__a21oi_1 _25188_ (.A1(_00914_),
    .A2(_00927_),
    .B1(_00926_),
    .Y(_00929_));
 sky130_fd_sc_hd__a31oi_2 _25189_ (.A1(_00551_),
    .A2(_00556_),
    .A3(_00559_),
    .B1(_00552_),
    .Y(_00930_));
 sky130_fd_sc_hd__a31o_1 _25190_ (.A1(_00551_),
    .A2(_00556_),
    .A3(_00559_),
    .B1(_00552_),
    .X(_00932_));
 sky130_fd_sc_hd__nand2_1 _25191_ (.A(_00932_),
    .B(_00929_),
    .Y(_00933_));
 sky130_fd_sc_hd__o21ai_1 _25192_ (.A1(_00926_),
    .A2(_00928_),
    .B1(_00930_),
    .Y(_00934_));
 sky130_fd_sc_hd__o311a_2 _25193_ (.A1(_00926_),
    .A2(_00928_),
    .A3(_00930_),
    .B1(net278),
    .C1(_00934_),
    .X(_00935_));
 sky130_fd_sc_hd__nor2_1 _25194_ (.A(_00925_),
    .B(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__o22a_2 _25195_ (.A1(_03986_),
    .A2(_03997_),
    .B1(_00925_),
    .B2(_00935_),
    .X(_00937_));
 sky130_fd_sc_hd__or3_2 _25196_ (.A(net302),
    .B(_04019_),
    .C(_00936_),
    .X(_00938_));
 sky130_fd_sc_hd__a311o_4 _25197_ (.A1(_00933_),
    .A2(_00934_),
    .A3(net278),
    .B1(net151),
    .C1(_00925_),
    .X(_00939_));
 sky130_fd_sc_hd__o22a_1 _25198_ (.A1(net170),
    .A2(net169),
    .B1(_00925_),
    .B2(_00935_),
    .X(_00940_));
 sky130_fd_sc_hd__o22ai_4 _25199_ (.A1(net170),
    .A2(net169),
    .B1(_00925_),
    .B2(_00935_),
    .Y(_00941_));
 sky130_fd_sc_hd__nand2_1 _25200_ (.A(_00939_),
    .B(_00941_),
    .Y(_00943_));
 sky130_fd_sc_hd__and3_1 _25201_ (.A(_14286_),
    .B(_14287_),
    .C(_13890_),
    .X(_00944_));
 sky130_fd_sc_hd__nand3_1 _25202_ (.A(_00570_),
    .B(_00944_),
    .C(_00213_),
    .Y(_00945_));
 sky130_fd_sc_hd__o211ai_4 _25203_ (.A1(_00568_),
    .A2(_00574_),
    .B1(_00945_),
    .C1(_00572_),
    .Y(_00946_));
 sky130_fd_sc_hd__nand4_1 _25204_ (.A(_00944_),
    .B(_00212_),
    .C(_00210_),
    .D(_13904_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand3b_4 _25205_ (.A_N(_00947_),
    .B(_00572_),
    .C(_00570_),
    .Y(_00948_));
 sky130_fd_sc_hd__nand2_1 _25206_ (.A(_00946_),
    .B(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__a22oi_1 _25207_ (.A1(_00939_),
    .A2(_00941_),
    .B1(_00946_),
    .B2(_00948_),
    .Y(_00950_));
 sky130_fd_sc_hd__a22o_2 _25208_ (.A1(_00939_),
    .A2(_00941_),
    .B1(_00946_),
    .B2(_00948_),
    .X(_00951_));
 sky130_fd_sc_hd__nand4_4 _25209_ (.A(_00939_),
    .B(_00941_),
    .C(_00946_),
    .D(_00948_),
    .Y(_00952_));
 sky130_fd_sc_hd__o22ai_1 _25210_ (.A1(net302),
    .A2(_04019_),
    .B1(_00943_),
    .B2(_00949_),
    .Y(_00954_));
 sky130_fd_sc_hd__nand3_2 _25211_ (.A(_00951_),
    .B(_00952_),
    .C(_04029_),
    .Y(_00955_));
 sky130_fd_sc_hd__a31oi_1 _25212_ (.A1(_00951_),
    .A2(_00952_),
    .A3(_04029_),
    .B1(_00937_),
    .Y(_00956_));
 sky130_fd_sc_hd__o22ai_2 _25213_ (.A1(_04029_),
    .A2(_00936_),
    .B1(_00950_),
    .B2(_00954_),
    .Y(_00957_));
 sky130_fd_sc_hd__a21oi_4 _25214_ (.A1(_00938_),
    .A2(_00955_),
    .B1(net271),
    .Y(_00958_));
 sky130_fd_sc_hd__or3_2 _25215_ (.A(net296),
    .B(_05232_),
    .C(_00956_),
    .X(_00959_));
 sky130_fd_sc_hd__a31o_1 _25216_ (.A1(_00951_),
    .A2(_00952_),
    .A3(_04029_),
    .B1(net171),
    .X(_00960_));
 sky130_fd_sc_hd__a311oi_4 _25217_ (.A1(_00951_),
    .A2(_00952_),
    .A3(_04029_),
    .B1(net171),
    .C1(_00937_),
    .Y(_00961_));
 sky130_fd_sc_hd__nand3_2 _25218_ (.A(_00955_),
    .B(net172),
    .C(_00938_),
    .Y(_00962_));
 sky130_fd_sc_hd__a2bb2oi_2 _25219_ (.A1_N(net189),
    .A2_N(net188),
    .B1(_00938_),
    .B2(_00955_),
    .Y(_00963_));
 sky130_fd_sc_hd__o21ai_4 _25220_ (.A1(net189),
    .A2(net188),
    .B1(_00957_),
    .Y(_00965_));
 sky130_fd_sc_hd__a31o_1 _25221_ (.A1(_00224_),
    .A2(_00581_),
    .A3(_00586_),
    .B1(_00587_),
    .X(_00966_));
 sky130_fd_sc_hd__o22ai_4 _25222_ (.A1(_00566_),
    .A2(_00584_),
    .B1(_00587_),
    .B2(_00583_),
    .Y(_00967_));
 sky130_fd_sc_hd__o21ai_4 _25223_ (.A1(_00961_),
    .A2(_00963_),
    .B1(_00967_),
    .Y(_00968_));
 sky130_fd_sc_hd__o211ai_4 _25224_ (.A1(_00937_),
    .A2(_00960_),
    .B1(_00966_),
    .C1(_00965_),
    .Y(_00969_));
 sky130_fd_sc_hd__o311a_1 _25225_ (.A1(_00961_),
    .A2(_00963_),
    .A3(_00967_),
    .B1(net271),
    .C1(_00968_),
    .X(_00970_));
 sky130_fd_sc_hd__nand3_4 _25226_ (.A(_00968_),
    .B(_00969_),
    .C(net271),
    .Y(_00971_));
 sky130_fd_sc_hd__o31a_1 _25227_ (.A1(net296),
    .A2(_05232_),
    .A3(_00956_),
    .B1(_00971_),
    .X(_00972_));
 sky130_fd_sc_hd__a31o_1 _25228_ (.A1(_00968_),
    .A2(_00969_),
    .A3(net271),
    .B1(_00958_),
    .X(_00973_));
 sky130_fd_sc_hd__o311a_1 _25229_ (.A1(_08311_),
    .A2(net215),
    .A3(_00235_),
    .B1(_00603_),
    .C1(_00608_),
    .X(_00974_));
 sky130_fd_sc_hd__o221ai_4 _25230_ (.A1(net200),
    .A2(_00235_),
    .B1(net177),
    .B2(_00598_),
    .C1(_00608_),
    .Y(_00976_));
 sky130_fd_sc_hd__a21oi_1 _25231_ (.A1(_00239_),
    .A2(_00608_),
    .B1(_00604_),
    .Y(_00977_));
 sky130_fd_sc_hd__a311oi_4 _25232_ (.A1(_00968_),
    .A2(_00969_),
    .A3(net271),
    .B1(net173),
    .C1(_00958_),
    .Y(_00978_));
 sky130_fd_sc_hd__nand3_4 _25233_ (.A(_00971_),
    .B(net174),
    .C(_00959_),
    .Y(_00979_));
 sky130_fd_sc_hd__a2bb2oi_4 _25234_ (.A1_N(_09134_),
    .A2_N(net192),
    .B1(_00959_),
    .B2(_00971_),
    .Y(_00980_));
 sky130_fd_sc_hd__o22ai_4 _25235_ (.A1(_09134_),
    .A2(net192),
    .B1(_00958_),
    .B2(_00970_),
    .Y(_00981_));
 sky130_fd_sc_hd__nor2_1 _25236_ (.A(_00978_),
    .B(_00980_),
    .Y(_00982_));
 sky130_fd_sc_hd__o211ai_1 _25237_ (.A1(_00604_),
    .A2(_00974_),
    .B1(_00979_),
    .C1(_00981_),
    .Y(_00983_));
 sky130_fd_sc_hd__o22ai_1 _25238_ (.A1(_00601_),
    .A2(_00977_),
    .B1(_00978_),
    .B2(_00980_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand3_1 _25239_ (.A(_00983_),
    .B(_00984_),
    .C(net244),
    .Y(_00985_));
 sky130_fd_sc_hd__a211o_1 _25240_ (.A1(_00959_),
    .A2(_00971_),
    .B1(net270),
    .C1(net268),
    .X(_00987_));
 sky130_fd_sc_hd__o2111ai_4 _25241_ (.A1(net175),
    .A2(_00599_),
    .B1(_00976_),
    .C1(_00979_),
    .D1(_00981_),
    .Y(_00988_));
 sky130_fd_sc_hd__o22ai_2 _25242_ (.A1(_00604_),
    .A2(_00974_),
    .B1(_00978_),
    .B2(_00980_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand3_4 _25243_ (.A(_00988_),
    .B(_00989_),
    .C(net244),
    .Y(_00990_));
 sky130_fd_sc_hd__o21ai_4 _25244_ (.A1(net244),
    .A2(_00972_),
    .B1(_00990_),
    .Y(_00991_));
 sky130_fd_sc_hd__inv_2 _25245_ (.A(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__o311a_2 _25246_ (.A1(net270),
    .A2(net268),
    .A3(_00972_),
    .B1(_00990_),
    .C1(_05754_),
    .X(_00993_));
 sky130_fd_sc_hd__o211ai_4 _25247_ (.A1(_00973_),
    .A2(net244),
    .B1(net175),
    .C1(_00985_),
    .Y(_00994_));
 sky130_fd_sc_hd__nand3_4 _25248_ (.A(_00990_),
    .B(net177),
    .C(_00987_),
    .Y(_00995_));
 sky130_fd_sc_hd__nand2_1 _25249_ (.A(_00994_),
    .B(_00995_),
    .Y(_00996_));
 sky130_fd_sc_hd__o21ai_2 _25250_ (.A1(net198),
    .A2(_00617_),
    .B1(_00634_),
    .Y(_00998_));
 sky130_fd_sc_hd__o221ai_4 _25251_ (.A1(_13520_),
    .A2(_00633_),
    .B1(_00617_),
    .B2(_08314_),
    .C1(_00632_),
    .Y(_00999_));
 sky130_fd_sc_hd__o22ai_2 _25252_ (.A1(net200),
    .A2(_00618_),
    .B1(_00998_),
    .B2(_00631_),
    .Y(_01000_));
 sky130_fd_sc_hd__o2111a_1 _25253_ (.A1(net200),
    .A2(_00618_),
    .B1(_00994_),
    .C1(_00995_),
    .D1(_00999_),
    .X(_01001_));
 sky130_fd_sc_hd__o2111ai_4 _25254_ (.A1(net199),
    .A2(_00618_),
    .B1(_00994_),
    .C1(_00995_),
    .D1(_00999_),
    .Y(_01002_));
 sky130_fd_sc_hd__a22o_2 _25255_ (.A1(_00994_),
    .A2(_00995_),
    .B1(_00999_),
    .B2(_00620_),
    .X(_01003_));
 sky130_fd_sc_hd__o2bb2ai_1 _25256_ (.A1_N(_00996_),
    .A2_N(_01000_),
    .B1(net265),
    .B2(net264),
    .Y(_01004_));
 sky130_fd_sc_hd__a211o_1 _25257_ (.A1(_00987_),
    .A2(_00990_),
    .B1(net265),
    .C1(net264),
    .X(_01005_));
 sky130_fd_sc_hd__nand3_1 _25258_ (.A(_01000_),
    .B(_00995_),
    .C(_00994_),
    .Y(_01006_));
 sky130_fd_sc_hd__o211ai_1 _25259_ (.A1(net200),
    .A2(_00618_),
    .B1(_00641_),
    .C1(_00996_),
    .Y(_01007_));
 sky130_fd_sc_hd__nand3_1 _25260_ (.A(_01006_),
    .B(_01007_),
    .C(net243),
    .Y(_01009_));
 sky130_fd_sc_hd__a31oi_4 _25261_ (.A1(_01003_),
    .A2(net243),
    .A3(_01002_),
    .B1(_00993_),
    .Y(_01010_));
 sky130_fd_sc_hd__a31o_4 _25262_ (.A1(_01003_),
    .A2(net243),
    .A3(_01002_),
    .B1(_00993_),
    .X(_01011_));
 sky130_fd_sc_hd__a311oi_4 _25263_ (.A1(_01003_),
    .A2(net243),
    .A3(_01002_),
    .B1(net200),
    .C1(_00993_),
    .Y(_01012_));
 sky130_fd_sc_hd__o221ai_4 _25264_ (.A1(net243),
    .A2(_00991_),
    .B1(_01001_),
    .B2(_01004_),
    .C1(net198),
    .Y(_01013_));
 sky130_fd_sc_hd__a31oi_1 _25265_ (.A1(_01006_),
    .A2(_01007_),
    .A3(net243),
    .B1(net198),
    .Y(_01014_));
 sky130_fd_sc_hd__nand3_2 _25266_ (.A(_01009_),
    .B(net200),
    .C(_01005_),
    .Y(_01015_));
 sky130_fd_sc_hd__a21oi_2 _25267_ (.A1(_01005_),
    .A2(_01014_),
    .B1(_01012_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_2 _25268_ (.A(_01013_),
    .B(_01015_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand4_2 _25269_ (.A(_13973_),
    .B(_13977_),
    .C(_14360_),
    .D(_14362_),
    .Y(_01018_));
 sky130_fd_sc_hd__a211oi_4 _25270_ (.A1(_00266_),
    .A2(_00281_),
    .B1(_01018_),
    .C1(_00285_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand2_1 _25271_ (.A(_00651_),
    .B(_01020_),
    .Y(_01021_));
 sky130_fd_sc_hd__a32oi_1 _25272_ (.A1(_00647_),
    .A2(_07934_),
    .A3(_07933_),
    .B1(_00651_),
    .B2(_01020_),
    .Y(_01022_));
 sky130_fd_sc_hd__o211a_2 _25273_ (.A1(_00656_),
    .A2(_00650_),
    .B1(_00652_),
    .C1(_01021_),
    .X(_01023_));
 sky130_fd_sc_hd__o211ai_4 _25274_ (.A1(_00656_),
    .A2(_00650_),
    .B1(_00652_),
    .C1(_01021_),
    .Y(_01024_));
 sky130_fd_sc_hd__o211ai_4 _25275_ (.A1(_13967_),
    .A2(_13970_),
    .B1(_01020_),
    .C1(_00652_),
    .Y(_01025_));
 sky130_fd_sc_hd__nand4_4 _25276_ (.A(_01020_),
    .B(_00652_),
    .C(_00651_),
    .D(_13971_),
    .Y(_01026_));
 sky130_fd_sc_hd__inv_2 _25277_ (.A(_01026_),
    .Y(_01027_));
 sky130_fd_sc_hd__a2bb2oi_1 _25278_ (.A1_N(_00650_),
    .A2_N(_01025_),
    .B1(_00661_),
    .B2(_01022_),
    .Y(_01028_));
 sky130_fd_sc_hd__o21ai_4 _25279_ (.A1(_00650_),
    .A2(_01025_),
    .B1(_01024_),
    .Y(_01029_));
 sky130_fd_sc_hd__a21oi_4 _25280_ (.A1(_01024_),
    .A2(_01026_),
    .B1(_01017_),
    .Y(_01031_));
 sky130_fd_sc_hd__a31o_2 _25281_ (.A1(_01017_),
    .A2(_01024_),
    .A3(_01026_),
    .B1(_05995_),
    .X(_01032_));
 sky130_fd_sc_hd__nand4_1 _25282_ (.A(_01013_),
    .B(_01015_),
    .C(_01024_),
    .D(_01026_),
    .Y(_01033_));
 sky130_fd_sc_hd__o221ai_4 _25283_ (.A1(net260),
    .A2(net255),
    .B1(_01016_),
    .B2(_01028_),
    .C1(_01033_),
    .Y(_01034_));
 sky130_fd_sc_hd__o221a_2 _25284_ (.A1(net240),
    .A2(_01010_),
    .B1(_01031_),
    .B2(_01032_),
    .C1(_06294_),
    .X(_01035_));
 sky130_fd_sc_hd__o221ai_4 _25285_ (.A1(net240),
    .A2(_01010_),
    .B1(_01031_),
    .B2(_01032_),
    .C1(_06294_),
    .Y(_01036_));
 sky130_fd_sc_hd__o311a_1 _25286_ (.A1(net260),
    .A2(net255),
    .A3(_01011_),
    .B1(_07935_),
    .C1(_01034_),
    .X(_01037_));
 sky130_fd_sc_hd__o211ai_4 _25287_ (.A1(net240),
    .A2(_01011_),
    .B1(_07935_),
    .C1(_01034_),
    .Y(_01038_));
 sky130_fd_sc_hd__o221ai_4 _25288_ (.A1(net240),
    .A2(_01010_),
    .B1(_01031_),
    .B2(_01032_),
    .C1(_07936_),
    .Y(_01039_));
 sky130_fd_sc_hd__a21oi_1 _25289_ (.A1(_00297_),
    .A2(_00666_),
    .B1(_00672_),
    .Y(_01040_));
 sky130_fd_sc_hd__a31o_1 _25290_ (.A1(_00297_),
    .A2(_00666_),
    .A3(_00671_),
    .B1(_00672_),
    .X(_01042_));
 sky130_fd_sc_hd__a31oi_4 _25291_ (.A1(_00297_),
    .A2(_00666_),
    .A3(_00671_),
    .B1(_00672_),
    .Y(_01043_));
 sky130_fd_sc_hd__o2bb2ai_4 _25292_ (.A1_N(_01038_),
    .A2_N(_01039_),
    .B1(_01040_),
    .B2(_00670_),
    .Y(_01044_));
 sky130_fd_sc_hd__nand3_4 _25293_ (.A(_01042_),
    .B(_01039_),
    .C(_01038_),
    .Y(_01045_));
 sky130_fd_sc_hd__nand3_2 _25294_ (.A(_01044_),
    .B(_01045_),
    .C(net214),
    .Y(_01046_));
 sky130_fd_sc_hd__a31oi_4 _25295_ (.A1(_01044_),
    .A2(_01045_),
    .A3(net214),
    .B1(_01035_),
    .Y(_01047_));
 sky130_fd_sc_hd__a311o_2 _25296_ (.A1(_01044_),
    .A2(_01045_),
    .A3(net214),
    .B1(net209),
    .C1(_01035_),
    .X(_01048_));
 sky130_fd_sc_hd__o211ai_4 _25297_ (.A1(_00308_),
    .A2(net227),
    .B1(_00685_),
    .C1(_00320_),
    .Y(_01049_));
 sky130_fd_sc_hd__o21ai_1 _25298_ (.A1(net223),
    .A2(_00683_),
    .B1(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__a311oi_4 _25299_ (.A1(_01044_),
    .A2(_01045_),
    .A3(net214),
    .B1(net202),
    .C1(_01035_),
    .Y(_01051_));
 sky130_fd_sc_hd__nand3_2 _25300_ (.A(_01046_),
    .B(_07564_),
    .C(_01036_),
    .Y(_01053_));
 sky130_fd_sc_hd__a2bb2oi_4 _25301_ (.A1_N(net221),
    .A2_N(net220),
    .B1(_01036_),
    .B2(_01046_),
    .Y(_01054_));
 sky130_fd_sc_hd__a22o_1 _25302_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_01036_),
    .B2(_01046_),
    .X(_01055_));
 sky130_fd_sc_hd__nand3_1 _25303_ (.A(_01050_),
    .B(_01053_),
    .C(_01055_),
    .Y(_01056_));
 sky130_fd_sc_hd__o221ai_4 _25304_ (.A1(net223),
    .A2(_00683_),
    .B1(_01051_),
    .B2(_01054_),
    .C1(_01049_),
    .Y(_01057_));
 sky130_fd_sc_hd__o211ai_4 _25305_ (.A1(net238),
    .A2(_06610_),
    .B1(_01056_),
    .C1(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__a21oi_1 _25306_ (.A1(_01036_),
    .A2(_01046_),
    .B1(net209),
    .Y(_01059_));
 sky130_fd_sc_hd__or3_1 _25307_ (.A(net238),
    .B(_06610_),
    .C(_01047_),
    .X(_01060_));
 sky130_fd_sc_hd__o2111ai_2 _25308_ (.A1(net223),
    .A2(_00683_),
    .B1(_01049_),
    .C1(_01053_),
    .D1(_01055_),
    .Y(_01061_));
 sky130_fd_sc_hd__o21ai_1 _25309_ (.A1(_01051_),
    .A2(_01054_),
    .B1(_01050_),
    .Y(_01062_));
 sky130_fd_sc_hd__nand3_2 _25310_ (.A(_01061_),
    .B(_01062_),
    .C(net209),
    .Y(_01064_));
 sky130_fd_sc_hd__a31o_2 _25311_ (.A1(_01061_),
    .A2(_01062_),
    .A3(net209),
    .B1(_01059_),
    .X(_01065_));
 sky130_fd_sc_hd__nand2_2 _25312_ (.A(_01048_),
    .B(_01058_),
    .Y(_01066_));
 sky130_fd_sc_hd__a2bb2oi_1 _25313_ (.A1_N(_07242_),
    .A2_N(net248),
    .B1(_01060_),
    .B2(_01064_),
    .Y(_01067_));
 sky130_fd_sc_hd__o211ai_4 _25314_ (.A1(_07242_),
    .A2(net248),
    .B1(_01048_),
    .C1(_01058_),
    .Y(_01068_));
 sky130_fd_sc_hd__o211a_1 _25315_ (.A1(net210),
    .A2(_01047_),
    .B1(_07246_),
    .C1(_01064_),
    .X(_01069_));
 sky130_fd_sc_hd__o211ai_4 _25316_ (.A1(net210),
    .A2(_01047_),
    .B1(_07246_),
    .C1(_01064_),
    .Y(_01070_));
 sky130_fd_sc_hd__nor2_1 _25317_ (.A(_01067_),
    .B(_01069_),
    .Y(_01071_));
 sky130_fd_sc_hd__nand2_1 _25318_ (.A(_01068_),
    .B(_01070_),
    .Y(_01072_));
 sky130_fd_sc_hd__a31oi_4 _25319_ (.A1(_00700_),
    .A2(_00706_),
    .A3(_00709_),
    .B1(_00697_),
    .Y(_01073_));
 sky130_fd_sc_hd__nand4_1 _25320_ (.A(_00698_),
    .B(_00715_),
    .C(_01068_),
    .D(_01070_),
    .Y(_01075_));
 sky130_fd_sc_hd__o221ai_4 _25321_ (.A1(net231),
    .A2(net228),
    .B1(_01073_),
    .B2(_01071_),
    .C1(_01075_),
    .Y(_01076_));
 sky130_fd_sc_hd__o221a_1 _25322_ (.A1(_06922_),
    .A2(_00694_),
    .B1(_01067_),
    .B2(_01069_),
    .C1(_00716_),
    .X(_01077_));
 sky130_fd_sc_hd__o22ai_2 _25323_ (.A1(net229),
    .A2(net228),
    .B1(_01072_),
    .B2(_01073_),
    .Y(_01078_));
 sky130_fd_sc_hd__o22a_2 _25324_ (.A1(net208),
    .A2(_01066_),
    .B1(_01077_),
    .B2(_01078_),
    .X(_01079_));
 sky130_fd_sc_hd__inv_2 _25325_ (.A(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__o211a_1 _25326_ (.A1(net208),
    .A2(_01065_),
    .B1(_01076_),
    .C1(_06924_),
    .X(_01081_));
 sky130_fd_sc_hd__o211ai_2 _25327_ (.A1(net208),
    .A2(_01065_),
    .B1(_01076_),
    .C1(_06924_),
    .Y(_01082_));
 sky130_fd_sc_hd__o221ai_4 _25328_ (.A1(net208),
    .A2(_01066_),
    .B1(_01077_),
    .B2(_01078_),
    .C1(_06922_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand2_1 _25329_ (.A(_01082_),
    .B(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hd__and4_1 _25330_ (.A(_14039_),
    .B(_14040_),
    .C(_14433_),
    .D(_14435_),
    .X(_01086_));
 sky130_fd_sc_hd__nand3_1 _25331_ (.A(_00724_),
    .B(_01086_),
    .C(_00353_),
    .Y(_01087_));
 sky130_fd_sc_hd__o211ai_4 _25332_ (.A1(_00728_),
    .A2(_00722_),
    .B1(_00725_),
    .C1(_01087_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand4_1 _25333_ (.A(_01086_),
    .B(_00352_),
    .C(_00349_),
    .D(_14048_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand3b_4 _25334_ (.A_N(_01089_),
    .B(_00725_),
    .C(_00724_),
    .Y(_01090_));
 sky130_fd_sc_hd__nand2_1 _25335_ (.A(_01088_),
    .B(_01090_),
    .Y(_01091_));
 sky130_fd_sc_hd__a21oi_2 _25336_ (.A1(_01088_),
    .A2(_01090_),
    .B1(_01084_),
    .Y(_01092_));
 sky130_fd_sc_hd__a21o_1 _25337_ (.A1(_01088_),
    .A2(_01090_),
    .B1(_01084_),
    .X(_01093_));
 sky130_fd_sc_hd__a31oi_1 _25338_ (.A1(_01084_),
    .A2(_01088_),
    .A3(_01090_),
    .B1(_07232_),
    .Y(_01094_));
 sky130_fd_sc_hd__a31o_1 _25339_ (.A1(_01084_),
    .A2(_01088_),
    .A3(_01090_),
    .B1(_07232_),
    .X(_01095_));
 sky130_fd_sc_hd__a22o_1 _25340_ (.A1(_01082_),
    .A2(_01083_),
    .B1(_01088_),
    .B2(_01090_),
    .X(_01097_));
 sky130_fd_sc_hd__nand3_4 _25341_ (.A(_01083_),
    .B(_01088_),
    .C(_01090_),
    .Y(_01098_));
 sky130_fd_sc_hd__or3_1 _25342_ (.A(net207),
    .B(net205),
    .C(_01079_),
    .X(_01099_));
 sky130_fd_sc_hd__o221ai_4 _25343_ (.A1(net207),
    .A2(net205),
    .B1(_01081_),
    .B2(_01098_),
    .C1(_01097_),
    .Y(_01100_));
 sky130_fd_sc_hd__a2bb2oi_1 _25344_ (.A1_N(_07233_),
    .A2_N(_01080_),
    .B1(_01093_),
    .B2(_01094_),
    .Y(_01101_));
 sky130_fd_sc_hd__a22o_1 _25345_ (.A1(_07232_),
    .A2(_01079_),
    .B1(_01094_),
    .B2(_01093_),
    .X(_01102_));
 sky130_fd_sc_hd__o221a_4 _25346_ (.A1(_07233_),
    .A2(_01080_),
    .B1(_01092_),
    .B2(_01095_),
    .C1(_07550_),
    .X(_01103_));
 sky130_fd_sc_hd__inv_2 _25347_ (.A(_01103_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand3_4 _25348_ (.A(_01100_),
    .B(net235),
    .C(_01099_),
    .Y(_01105_));
 sky130_fd_sc_hd__o221ai_4 _25349_ (.A1(_07233_),
    .A2(_01080_),
    .B1(_01092_),
    .B2(_01095_),
    .C1(net233),
    .Y(_01106_));
 sky130_fd_sc_hd__o21a_1 _25350_ (.A1(_00365_),
    .A2(_00739_),
    .B1(_00748_),
    .X(_01108_));
 sky130_fd_sc_hd__a21oi_1 _25351_ (.A1(_00364_),
    .A2(_00740_),
    .B1(_00746_),
    .Y(_01109_));
 sky130_fd_sc_hd__o21ai_2 _25352_ (.A1(_00746_),
    .A2(_00742_),
    .B1(_00748_),
    .Y(_01110_));
 sky130_fd_sc_hd__a21oi_1 _25353_ (.A1(_01105_),
    .A2(_01106_),
    .B1(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__o2bb2ai_2 _25354_ (.A1_N(_01105_),
    .A2_N(_01106_),
    .B1(_01108_),
    .B2(_00746_),
    .Y(_01112_));
 sky130_fd_sc_hd__o211a_1 _25355_ (.A1(_00747_),
    .A2(_01109_),
    .B1(_01106_),
    .C1(_01105_),
    .X(_01113_));
 sky130_fd_sc_hd__nand3_4 _25356_ (.A(_01105_),
    .B(_01106_),
    .C(_01110_),
    .Y(_01114_));
 sky130_fd_sc_hd__o21ai_1 _25357_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_01114_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand3_1 _25358_ (.A(_01112_),
    .B(_01114_),
    .C(net163),
    .Y(_01116_));
 sky130_fd_sc_hd__or3_1 _25359_ (.A(_07544_),
    .B(_07546_),
    .C(_01101_),
    .X(_01117_));
 sky130_fd_sc_hd__o22ai_2 _25360_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_01111_),
    .B2(_01113_),
    .Y(_01119_));
 sky130_fd_sc_hd__a31o_1 _25361_ (.A1(_01112_),
    .A2(_01114_),
    .A3(net163),
    .B1(_01103_),
    .X(_01120_));
 sky130_fd_sc_hd__o211a_1 _25362_ (.A1(_00386_),
    .A2(_00381_),
    .B1(_00379_),
    .C1(_00760_),
    .X(_01121_));
 sky130_fd_sc_hd__and3_1 _25363_ (.A(_00382_),
    .B(_00762_),
    .C(_00764_),
    .X(_01122_));
 sky130_fd_sc_hd__a31o_1 _25364_ (.A1(_00382_),
    .A2(_00762_),
    .A3(_00764_),
    .B1(_00759_),
    .X(_01123_));
 sky130_fd_sc_hd__o21ai_2 _25365_ (.A1(_01111_),
    .A2(_01115_),
    .B1(_06314_),
    .Y(_01124_));
 sky130_fd_sc_hd__a311oi_2 _25366_ (.A1(_01112_),
    .A2(_01114_),
    .A3(net163),
    .B1(_01103_),
    .C1(net252),
    .Y(_01125_));
 sky130_fd_sc_hd__a311o_1 _25367_ (.A1(_01112_),
    .A2(_01114_),
    .A3(net163),
    .B1(_01103_),
    .C1(net252),
    .X(_01126_));
 sky130_fd_sc_hd__a2bb2oi_2 _25368_ (.A1_N(net284),
    .A2_N(net281),
    .B1(_01104_),
    .B2(_01116_),
    .Y(_01127_));
 sky130_fd_sc_hd__o211ai_4 _25369_ (.A1(net284),
    .A2(net282),
    .B1(_01117_),
    .C1(_01119_),
    .Y(_01128_));
 sky130_fd_sc_hd__o221ai_2 _25370_ (.A1(_00761_),
    .A2(_01121_),
    .B1(_01103_),
    .B2(_01124_),
    .C1(_01128_),
    .Y(_01130_));
 sky130_fd_sc_hd__o22ai_1 _25371_ (.A1(_00759_),
    .A2(_01122_),
    .B1(_01125_),
    .B2(_01127_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand3_2 _25372_ (.A(_01131_),
    .B(net162),
    .C(_01130_),
    .Y(_01132_));
 sky130_fd_sc_hd__a211o_2 _25373_ (.A1(_01104_),
    .A2(_01116_),
    .B1(net183),
    .C1(net182),
    .X(_01133_));
 sky130_fd_sc_hd__o211ai_2 _25374_ (.A1(_01103_),
    .A2(_01124_),
    .B1(_01123_),
    .C1(_01128_),
    .Y(_01134_));
 sky130_fd_sc_hd__o22ai_2 _25375_ (.A1(_00761_),
    .A2(_01121_),
    .B1(_01125_),
    .B2(_01127_),
    .Y(_01135_));
 sky130_fd_sc_hd__o211ai_4 _25376_ (.A1(net183),
    .A2(net182),
    .B1(_01134_),
    .C1(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__o21a_2 _25377_ (.A1(net162),
    .A2(_01120_),
    .B1(_01132_),
    .X(_01137_));
 sky130_fd_sc_hd__and3_1 _25378_ (.A(_08301_),
    .B(_01133_),
    .C(_01136_),
    .X(_01138_));
 sky130_fd_sc_hd__a2bb2oi_4 _25379_ (.A1_N(_06009_),
    .A2_N(net287),
    .B1(_01133_),
    .B2(_01136_),
    .Y(_01139_));
 sky130_fd_sc_hd__o211ai_4 _25380_ (.A1(_01120_),
    .A2(net162),
    .B1(_06014_),
    .C1(_01132_),
    .Y(_01141_));
 sky130_fd_sc_hd__o211a_2 _25381_ (.A1(net285),
    .A2(_06012_),
    .B1(_01133_),
    .C1(_01136_),
    .X(_01142_));
 sky130_fd_sc_hd__o211ai_4 _25382_ (.A1(net285),
    .A2(_06012_),
    .B1(_01133_),
    .C1(_01136_),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_1 _25383_ (.A(_01139_),
    .B(_01142_),
    .Y(_01144_));
 sky130_fd_sc_hd__o22ai_2 _25384_ (.A1(net263),
    .A2(_00771_),
    .B1(_00796_),
    .B2(_00785_),
    .Y(_01145_));
 sky130_fd_sc_hd__a31oi_1 _25385_ (.A1(_00779_),
    .A2(_00786_),
    .A3(_00790_),
    .B1(_00774_),
    .Y(_01146_));
 sky130_fd_sc_hd__nand4_4 _25386_ (.A(_00775_),
    .B(_00797_),
    .C(_01141_),
    .D(_01143_),
    .Y(_01147_));
 sky130_fd_sc_hd__o2bb2ai_4 _25387_ (.A1_N(_00775_),
    .A2_N(_00797_),
    .B1(_01139_),
    .B2(_01142_),
    .Y(_01148_));
 sky130_fd_sc_hd__o211ai_2 _25388_ (.A1(_08296_),
    .A2(net179),
    .B1(_01147_),
    .C1(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__and3_1 _25389_ (.A(_01137_),
    .B(_08299_),
    .C(_08297_),
    .X(_01150_));
 sky130_fd_sc_hd__a211o_1 _25390_ (.A1(_01133_),
    .A2(_01136_),
    .B1(_08296_),
    .C1(net179),
    .X(_01152_));
 sky130_fd_sc_hd__o21ai_2 _25391_ (.A1(_01139_),
    .A2(_01142_),
    .B1(_01146_),
    .Y(_01153_));
 sky130_fd_sc_hd__nand3_2 _25392_ (.A(_01145_),
    .B(_01143_),
    .C(_01141_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand3_1 _25393_ (.A(_01153_),
    .B(_01154_),
    .C(net159),
    .Y(_01155_));
 sky130_fd_sc_hd__a31o_1 _25394_ (.A1(_01148_),
    .A2(net159),
    .A3(_01147_),
    .B1(_01138_),
    .X(_01156_));
 sky130_fd_sc_hd__a311o_1 _25395_ (.A1(_01153_),
    .A2(_01154_),
    .A3(net159),
    .B1(net149),
    .C1(_01150_),
    .X(_01157_));
 sky130_fd_sc_hd__a311oi_4 _25396_ (.A1(_01148_),
    .A2(net159),
    .A3(_01147_),
    .B1(_01138_),
    .C1(net263),
    .Y(_01158_));
 sky130_fd_sc_hd__o211ai_4 _25397_ (.A1(net159),
    .A2(_01137_),
    .B1(_01149_),
    .C1(_05768_),
    .Y(_01159_));
 sky130_fd_sc_hd__a311oi_4 _25398_ (.A1(_01153_),
    .A2(_01154_),
    .A3(net159),
    .B1(_01150_),
    .C1(_05768_),
    .Y(_01160_));
 sky130_fd_sc_hd__nand3_4 _25399_ (.A(_01155_),
    .B(net263),
    .C(_01152_),
    .Y(_01161_));
 sky130_fd_sc_hd__o21ai_1 _25400_ (.A1(_05507_),
    .A2(_00802_),
    .B1(_00812_),
    .Y(_01163_));
 sky130_fd_sc_hd__o22ai_4 _25401_ (.A1(_00805_),
    .A2(_00772_),
    .B1(_00810_),
    .B2(_00808_),
    .Y(_01164_));
 sky130_fd_sc_hd__o211ai_4 _25402_ (.A1(_00808_),
    .A2(_00810_),
    .B1(_01161_),
    .C1(_00807_),
    .Y(_01165_));
 sky130_fd_sc_hd__nand4_2 _25403_ (.A(_00807_),
    .B(_01159_),
    .C(_01161_),
    .D(_01163_),
    .Y(_01166_));
 sky130_fd_sc_hd__o21ai_4 _25404_ (.A1(_01158_),
    .A2(_01160_),
    .B1(_01164_),
    .Y(_01167_));
 sky130_fd_sc_hd__nand3_1 _25405_ (.A(_01159_),
    .B(_01161_),
    .C(_01164_),
    .Y(_01168_));
 sky130_fd_sc_hd__o221ai_2 _25406_ (.A1(_00808_),
    .A2(_00810_),
    .B1(_01158_),
    .B2(_01160_),
    .C1(_00807_),
    .Y(_01169_));
 sky130_fd_sc_hd__o211ai_2 _25407_ (.A1(_08709_),
    .A2(_08712_),
    .B1(_01168_),
    .C1(_01169_),
    .Y(_01170_));
 sky130_fd_sc_hd__o211a_1 _25408_ (.A1(net159),
    .A2(_01137_),
    .B1(_01149_),
    .C1(_08715_),
    .X(_01171_));
 sky130_fd_sc_hd__a311o_2 _25409_ (.A1(_01148_),
    .A2(net159),
    .A3(_01147_),
    .B1(net149),
    .C1(_01138_),
    .X(_01172_));
 sky130_fd_sc_hd__o221ai_4 _25410_ (.A1(_08709_),
    .A2(_08712_),
    .B1(_01158_),
    .B2(_01165_),
    .C1(_01167_),
    .Y(_01174_));
 sky130_fd_sc_hd__a31o_1 _25411_ (.A1(_01167_),
    .A2(net149),
    .A3(_01166_),
    .B1(_01171_),
    .X(_01175_));
 sky130_fd_sc_hd__o21ai_2 _25412_ (.A1(_05248_),
    .A2(_00819_),
    .B1(_00825_),
    .Y(_01176_));
 sky130_fd_sc_hd__a21oi_1 _25413_ (.A1(_00827_),
    .A2(_00824_),
    .B1(_00828_),
    .Y(_01177_));
 sky130_fd_sc_hd__a311oi_4 _25414_ (.A1(_01167_),
    .A2(net149),
    .A3(_01166_),
    .B1(_01171_),
    .C1(net292),
    .Y(_01178_));
 sky130_fd_sc_hd__nand3_4 _25415_ (.A(_01174_),
    .B(_05507_),
    .C(_01172_),
    .Y(_01179_));
 sky130_fd_sc_hd__a22oi_1 _25416_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_01172_),
    .B2(_01174_),
    .Y(_01180_));
 sky130_fd_sc_hd__o211ai_4 _25417_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_01157_),
    .C1(_01170_),
    .Y(_01181_));
 sky130_fd_sc_hd__o2111a_1 _25418_ (.A1(_05249_),
    .A2(_00820_),
    .B1(_01176_),
    .C1(_01179_),
    .D1(_01181_),
    .X(_01182_));
 sky130_fd_sc_hd__o2111ai_4 _25419_ (.A1(_05249_),
    .A2(_00820_),
    .B1(_01176_),
    .C1(_01179_),
    .D1(_01181_),
    .Y(_01183_));
 sky130_fd_sc_hd__a22oi_1 _25420_ (.A1(_00827_),
    .A2(_01176_),
    .B1(_01179_),
    .B2(_01181_),
    .Y(_01185_));
 sky130_fd_sc_hd__o2bb2ai_1 _25421_ (.A1_N(_00827_),
    .A2_N(_01176_),
    .B1(_01178_),
    .B2(_01180_),
    .Y(_01186_));
 sky130_fd_sc_hd__o22ai_2 _25422_ (.A1(_09120_),
    .A2(net147),
    .B1(_01182_),
    .B2(_01185_),
    .Y(_01187_));
 sky130_fd_sc_hd__a211o_1 _25423_ (.A1(_01172_),
    .A2(_01174_),
    .B1(_09120_),
    .C1(net147),
    .X(_01188_));
 sky130_fd_sc_hd__o211ai_4 _25424_ (.A1(_09120_),
    .A2(net147),
    .B1(_01183_),
    .C1(_01186_),
    .Y(_01189_));
 sky130_fd_sc_hd__a211o_2 _25425_ (.A1(_01188_),
    .A2(_01189_),
    .B1(_09553_),
    .C1(net155),
    .X(_01190_));
 sky130_fd_sc_hd__inv_2 _25426_ (.A(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__a2bb2oi_2 _25427_ (.A1_N(net318),
    .A2_N(net315),
    .B1(_01188_),
    .B2(_01189_),
    .Y(_01192_));
 sky130_fd_sc_hd__o221ai_4 _25428_ (.A1(net318),
    .A2(net315),
    .B1(net146),
    .B2(_01175_),
    .C1(_01187_),
    .Y(_01193_));
 sky130_fd_sc_hd__o211a_2 _25429_ (.A1(_05246_),
    .A2(_05247_),
    .B1(_01188_),
    .C1(_01189_),
    .X(_01194_));
 sky130_fd_sc_hd__o211ai_1 _25430_ (.A1(_05246_),
    .A2(_05247_),
    .B1(_01188_),
    .C1(_01189_),
    .Y(_01196_));
 sky130_fd_sc_hd__o2bb2ai_4 _25431_ (.A1_N(_00840_),
    .A2_N(_00845_),
    .B1(_00841_),
    .B2(_00834_),
    .Y(_01197_));
 sky130_fd_sc_hd__o21ai_2 _25432_ (.A1(_01192_),
    .A2(_01194_),
    .B1(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__o311a_1 _25433_ (.A1(_01192_),
    .A2(_01197_),
    .A3(_01194_),
    .B1(net143),
    .C1(_01198_),
    .X(_01199_));
 sky130_fd_sc_hd__o311ai_4 _25434_ (.A1(_01192_),
    .A2(_01197_),
    .A3(_01194_),
    .B1(net143),
    .C1(_01198_),
    .Y(_01200_));
 sky130_fd_sc_hd__a2bb2oi_1 _25435_ (.A1_N(net340),
    .A2_N(_04184_),
    .B1(_01190_),
    .B2(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__o21ai_4 _25436_ (.A1(_01191_),
    .A2(_01199_),
    .B1(_04238_),
    .Y(_01202_));
 sky130_fd_sc_hd__o211a_1 _25437_ (.A1(_04206_),
    .A2(_04216_),
    .B1(_01190_),
    .C1(_01200_),
    .X(_01203_));
 sky130_fd_sc_hd__o211ai_4 _25438_ (.A1(_04206_),
    .A2(_04216_),
    .B1(_01190_),
    .C1(_01200_),
    .Y(_01204_));
 sky130_fd_sc_hd__a32o_1 _25439_ (.A1(_02104_),
    .A2(_02126_),
    .A3(_00851_),
    .B1(_00860_),
    .B2(_00861_),
    .X(_01205_));
 sky130_fd_sc_hd__a31oi_4 _25440_ (.A1(_00854_),
    .A2(_00860_),
    .A3(_00861_),
    .B1(_00852_),
    .Y(_01207_));
 sky130_fd_sc_hd__o21ai_2 _25441_ (.A1(_01201_),
    .A2(_01203_),
    .B1(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__o2111ai_4 _25442_ (.A1(_00851_),
    .A2(_02148_),
    .B1(_01204_),
    .C1(_01202_),
    .D1(_01205_),
    .Y(_01209_));
 sky130_fd_sc_hd__a22o_4 _25443_ (.A1(_09575_),
    .A2(_09577_),
    .B1(_01190_),
    .B2(_01200_),
    .X(_01210_));
 sky130_fd_sc_hd__o211ai_4 _25444_ (.A1(_09571_),
    .A2(_09573_),
    .B1(_01208_),
    .C1(_01209_),
    .Y(_01211_));
 sky130_fd_sc_hd__nand2_4 _25445_ (.A(_01210_),
    .B(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__a2bb2oi_4 _25446_ (.A1_N(_02049_),
    .A2_N(net343),
    .B1(_01210_),
    .B2(_01211_),
    .Y(_01213_));
 sky130_fd_sc_hd__a22o_4 _25447_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_01210_),
    .B2(_01211_),
    .X(_01214_));
 sky130_fd_sc_hd__a31oi_1 _25448_ (.A1(_09579_),
    .A2(_01208_),
    .A3(_01209_),
    .B1(_02148_),
    .Y(_01215_));
 sky130_fd_sc_hd__and3_2 _25449_ (.A(_01211_),
    .B(_02137_),
    .C(_01210_),
    .X(_01216_));
 sky130_fd_sc_hd__nand2_1 _25450_ (.A(_01215_),
    .B(_01210_),
    .Y(_01218_));
 sky130_fd_sc_hd__a21oi_1 _25451_ (.A1(_01210_),
    .A2(_01215_),
    .B1(_01213_),
    .Y(_01219_));
 sky130_fd_sc_hd__o2111ai_2 _25452_ (.A1(_14176_),
    .A2(_14167_),
    .B1(_14175_),
    .C1(_00112_),
    .D1(_00114_),
    .Y(_01220_));
 sky130_fd_sc_hd__nor3_1 _25453_ (.A(_00485_),
    .B(_01220_),
    .C(_00487_),
    .Y(_01221_));
 sky130_fd_sc_hd__nand2_1 _25454_ (.A(_01221_),
    .B(_00873_),
    .Y(_01222_));
 sky130_fd_sc_hd__o211ai_4 _25455_ (.A1(_00876_),
    .A2(_00872_),
    .B1(_00875_),
    .C1(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__nor4_1 _25456_ (.A(_14179_),
    .B(_00485_),
    .C(_01220_),
    .D(_00487_),
    .Y(_01224_));
 sky130_fd_sc_hd__nand3_4 _25457_ (.A(_00873_),
    .B(_00875_),
    .C(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_4 _25458_ (.A(_01223_),
    .B(_01225_),
    .Y(_01226_));
 sky130_fd_sc_hd__inv_2 _25459_ (.A(_01226_),
    .Y(_01227_));
 sky130_fd_sc_hd__o211a_1 _25460_ (.A1(_01213_),
    .A2(_01216_),
    .B1(_01223_),
    .C1(_01225_),
    .X(_01229_));
 sky130_fd_sc_hd__o2bb2ai_2 _25461_ (.A1_N(_01219_),
    .A2_N(_01226_),
    .B1(_10474_),
    .B2(net138),
    .Y(_01230_));
 sky130_fd_sc_hd__a21oi_1 _25462_ (.A1(_01210_),
    .A2(_01211_),
    .B1(net131),
    .Y(_01231_));
 sky130_fd_sc_hd__a211o_1 _25463_ (.A1(_01210_),
    .A2(_01211_),
    .B1(_10474_),
    .C1(net138),
    .X(_01232_));
 sky130_fd_sc_hd__o21ai_2 _25464_ (.A1(_01213_),
    .A2(_01216_),
    .B1(_01226_),
    .Y(_01233_));
 sky130_fd_sc_hd__o211ai_4 _25465_ (.A1(_02148_),
    .A2(_01212_),
    .B1(_01223_),
    .C1(_01225_),
    .Y(_01234_));
 sky130_fd_sc_hd__o2111ai_4 _25466_ (.A1(_01212_),
    .A2(_02148_),
    .B1(_01223_),
    .C1(_01214_),
    .D1(_01225_),
    .Y(_01235_));
 sky130_fd_sc_hd__o221ai_4 _25467_ (.A1(_10474_),
    .A2(net138),
    .B1(_01213_),
    .B2(_01234_),
    .C1(_01233_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor2_1 _25468_ (.A(_00885_),
    .B(_00891_),
    .Y(_01237_));
 sky130_fd_sc_hd__a311oi_4 _25469_ (.A1(net131),
    .A2(_01233_),
    .A3(_01235_),
    .B1(_01231_),
    .C1(_00251_),
    .Y(_01238_));
 sky130_fd_sc_hd__o211ai_2 _25470_ (.A1(_00218_),
    .A2(_00229_),
    .B1(_01232_),
    .C1(_01236_),
    .Y(_01240_));
 sky130_fd_sc_hd__o221a_1 _25471_ (.A1(net131),
    .A2(_01212_),
    .B1(_01229_),
    .B2(_01230_),
    .C1(_00251_),
    .X(_01241_));
 sky130_fd_sc_hd__o221ai_4 _25472_ (.A1(net131),
    .A2(_01212_),
    .B1(_01229_),
    .B2(_01230_),
    .C1(_00251_),
    .Y(_01242_));
 sky130_fd_sc_hd__o21ai_1 _25473_ (.A1(_00885_),
    .A2(_00891_),
    .B1(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__o21ai_1 _25474_ (.A1(_01238_),
    .A2(_01241_),
    .B1(_01237_),
    .Y(_01244_));
 sky130_fd_sc_hd__a211o_2 _25475_ (.A1(_01232_),
    .A2(_01236_),
    .B1(_10949_),
    .C1(net136),
    .X(_01245_));
 sky130_fd_sc_hd__o221ai_4 _25476_ (.A1(_10949_),
    .A2(net136),
    .B1(_01238_),
    .B2(_01243_),
    .C1(_01244_),
    .Y(_01246_));
 sky130_fd_sc_hd__nand2_1 _25477_ (.A(_01245_),
    .B(_01246_),
    .Y(_01247_));
 sky130_fd_sc_hd__a211o_1 _25478_ (.A1(_01245_),
    .A2(_01246_),
    .B1(_11459_),
    .C1(_11461_),
    .X(_01248_));
 sky130_fd_sc_hd__a21oi_1 _25479_ (.A1(_01245_),
    .A2(_01246_),
    .B1(_12888_),
    .Y(_01249_));
 sky130_fd_sc_hd__a211o_1 _25480_ (.A1(_01245_),
    .A2(_01246_),
    .B1(_12867_),
    .C1(_12877_),
    .X(_01251_));
 sky130_fd_sc_hd__and3_1 _25481_ (.A(_01246_),
    .B(_12888_),
    .C(_01245_),
    .X(_01252_));
 sky130_fd_sc_hd__o211ai_2 _25482_ (.A1(_12867_),
    .A2(_12877_),
    .B1(_01245_),
    .C1(_01246_),
    .Y(_01253_));
 sky130_fd_sc_hd__o21ai_1 _25483_ (.A1(_00895_),
    .A2(_00896_),
    .B1(_00898_),
    .Y(_01254_));
 sky130_fd_sc_hd__o221a_1 _25484_ (.A1(_00895_),
    .A2(_00896_),
    .B1(_01249_),
    .B2(_01252_),
    .C1(_00898_),
    .X(_01255_));
 sky130_fd_sc_hd__a31o_1 _25485_ (.A1(_01251_),
    .A2(_01253_),
    .A3(_01254_),
    .B1(_11464_),
    .X(_01256_));
 sky130_fd_sc_hd__a2bb2o_1 _25486_ (.A1_N(_01255_),
    .A2_N(_01256_),
    .B1(_11464_),
    .B2(_01247_),
    .X(_01257_));
 sky130_fd_sc_hd__and3_1 _25487_ (.A(_11265_),
    .B(_11287_),
    .C(_01257_),
    .X(_01258_));
 sky130_fd_sc_hd__o21ai_1 _25488_ (.A1(_11210_),
    .A2(_11232_),
    .B1(_01257_),
    .Y(_01259_));
 sky130_fd_sc_hd__o211a_1 _25489_ (.A1(_01255_),
    .A2(_01256_),
    .B1(_11298_),
    .C1(_01248_),
    .X(_01260_));
 sky130_fd_sc_hd__o32ai_4 _25490_ (.A1(_09927_),
    .A2(_09949_),
    .A3(_00903_),
    .B1(_00904_),
    .B2(_00906_),
    .Y(_01262_));
 sky130_fd_sc_hd__o21ai_1 _25491_ (.A1(_01258_),
    .A2(_01260_),
    .B1(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__a21o_1 _25492_ (.A1(_01263_),
    .A2(_11943_),
    .B1(_01257_),
    .X(_01264_));
 sky130_fd_sc_hd__xnor2_1 _25493_ (.A(_00912_),
    .B(_01264_),
    .Y(net99));
 sky130_fd_sc_hd__o31a_1 _25494_ (.A1(_00908_),
    .A2(_01264_),
    .A3(_00521_),
    .B1(_05119_),
    .X(_01265_));
 sky130_fd_sc_hd__a31o_1 _25495_ (.A1(_11471_),
    .A2(_00916_),
    .A3(_00921_),
    .B1(_00066_),
    .X(_01266_));
 sky130_fd_sc_hd__a311o_1 _25496_ (.A1(_11471_),
    .A2(_00916_),
    .A3(_00921_),
    .B1(net278),
    .C1(_00066_),
    .X(_01267_));
 sky130_fd_sc_hd__a21oi_1 _25497_ (.A1(_10963_),
    .A2(_10964_),
    .B1(_01266_),
    .Y(_01268_));
 sky130_fd_sc_hd__o21a_1 _25498_ (.A1(_10965_),
    .A2(_10967_),
    .B1(_01266_),
    .X(_01269_));
 sky130_fd_sc_hd__nor2_1 _25499_ (.A(_01268_),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__o21bai_1 _25500_ (.A1(_00928_),
    .A2(_00930_),
    .B1_N(_00926_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_1 _25501_ (.A(_01272_),
    .B(_01270_),
    .Y(_01273_));
 sky130_fd_sc_hd__o221ai_2 _25502_ (.A1(net150),
    .A2(_00924_),
    .B1(_01268_),
    .B2(_01269_),
    .C1(_00933_),
    .Y(_01274_));
 sky130_fd_sc_hd__nand3_1 _25503_ (.A(_01273_),
    .B(_01274_),
    .C(net278),
    .Y(_01275_));
 sky130_fd_sc_hd__o21a_2 _25504_ (.A1(net278),
    .A2(_01266_),
    .B1(_01275_),
    .X(_01276_));
 sky130_fd_sc_hd__or3_1 _25505_ (.A(net302),
    .B(_04019_),
    .C(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__a2bb2oi_1 _25506_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_01267_),
    .B2(_01275_),
    .Y(_01278_));
 sky130_fd_sc_hd__a2bb2o_1 _25507_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_01267_),
    .B2(_01275_),
    .X(_01279_));
 sky130_fd_sc_hd__a31oi_1 _25508_ (.A1(_01273_),
    .A2(_01274_),
    .A3(net278),
    .B1(_10492_),
    .Y(_01280_));
 sky130_fd_sc_hd__and3_1 _25509_ (.A(_01275_),
    .B(net150),
    .C(_01267_),
    .X(_01281_));
 sky130_fd_sc_hd__o21ai_1 _25510_ (.A1(net278),
    .A2(_01266_),
    .B1(_01280_),
    .Y(_01283_));
 sky130_fd_sc_hd__a21oi_1 _25511_ (.A1(_01267_),
    .A2(_01280_),
    .B1(_01278_),
    .Y(_01284_));
 sky130_fd_sc_hd__nand2_1 _25512_ (.A(_01279_),
    .B(_01283_),
    .Y(_01285_));
 sky130_fd_sc_hd__a31oi_4 _25513_ (.A1(_00939_),
    .A2(_00946_),
    .A3(_00948_),
    .B1(_00940_),
    .Y(_01286_));
 sky130_fd_sc_hd__a31o_1 _25514_ (.A1(_00939_),
    .A2(_00946_),
    .A3(_00948_),
    .B1(_00940_),
    .X(_01287_));
 sky130_fd_sc_hd__nand2_1 _25515_ (.A(_01287_),
    .B(_01284_),
    .Y(_01288_));
 sky130_fd_sc_hd__o221a_2 _25516_ (.A1(net153),
    .A2(_00936_),
    .B1(_01278_),
    .B2(_01281_),
    .C1(_00952_),
    .X(_01289_));
 sky130_fd_sc_hd__o21ai_1 _25517_ (.A1(_01278_),
    .A2(_01281_),
    .B1(_01286_),
    .Y(_01290_));
 sky130_fd_sc_hd__o22ai_4 _25518_ (.A1(net302),
    .A2(_04019_),
    .B1(_01286_),
    .B2(_01285_),
    .Y(_01291_));
 sky130_fd_sc_hd__nand3_1 _25519_ (.A(_01288_),
    .B(_01290_),
    .C(_04029_),
    .Y(_01292_));
 sky130_fd_sc_hd__o22ai_4 _25520_ (.A1(_04029_),
    .A2(_01276_),
    .B1(_01289_),
    .B2(_01291_),
    .Y(_01294_));
 sky130_fd_sc_hd__a211o_2 _25521_ (.A1(_01277_),
    .A2(_01292_),
    .B1(net296),
    .C1(_05232_),
    .X(_01295_));
 sky130_fd_sc_hd__inv_2 _25522_ (.A(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__a2bb2oi_1 _25523_ (.A1_N(net170),
    .A2_N(_10022_),
    .B1(_01277_),
    .B2(_01292_),
    .Y(_01297_));
 sky130_fd_sc_hd__o21ai_1 _25524_ (.A1(net170),
    .A2(_10022_),
    .B1(_01294_),
    .Y(_01298_));
 sky130_fd_sc_hd__o22a_1 _25525_ (.A1(net167),
    .A2(_10024_),
    .B1(_01289_),
    .B2(_01291_),
    .X(_01299_));
 sky130_fd_sc_hd__o221ai_4 _25526_ (.A1(_04029_),
    .A2(_01276_),
    .B1(_01289_),
    .B2(_01291_),
    .C1(net153),
    .Y(_01300_));
 sky130_fd_sc_hd__a21oi_1 _25527_ (.A1(_01299_),
    .A2(_01277_),
    .B1(_01297_),
    .Y(_01301_));
 sky130_fd_sc_hd__nand2_1 _25528_ (.A(_01298_),
    .B(_01300_),
    .Y(_01302_));
 sky130_fd_sc_hd__and4_1 _25529_ (.A(_14313_),
    .B(_14316_),
    .C(_00222_),
    .D(_00224_),
    .X(_01303_));
 sky130_fd_sc_hd__nand4_1 _25530_ (.A(_14313_),
    .B(_14316_),
    .C(_00222_),
    .D(_00224_),
    .Y(_01305_));
 sky130_fd_sc_hd__nor3_1 _25531_ (.A(_00585_),
    .B(_00587_),
    .C(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__nand3_1 _25532_ (.A(_00962_),
    .B(_01303_),
    .C(_00589_),
    .Y(_01307_));
 sky130_fd_sc_hd__o211ai_4 _25533_ (.A1(_00967_),
    .A2(_00961_),
    .B1(_00965_),
    .C1(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__nand4_4 _25534_ (.A(_01306_),
    .B(_00965_),
    .C(_00962_),
    .D(_14311_),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _25535_ (.A(_01308_),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__nand3_1 _25536_ (.A(_01302_),
    .B(_01308_),
    .C(_01309_),
    .Y(_01311_));
 sky130_fd_sc_hd__nand2_1 _25537_ (.A(_01310_),
    .B(_01301_),
    .Y(_01312_));
 sky130_fd_sc_hd__nand4_2 _25538_ (.A(_01298_),
    .B(_01300_),
    .C(_01308_),
    .D(_01309_),
    .Y(_01313_));
 sky130_fd_sc_hd__a22o_1 _25539_ (.A1(_01298_),
    .A2(_01300_),
    .B1(_01308_),
    .B2(_01309_),
    .X(_01314_));
 sky130_fd_sc_hd__nand3_2 _25540_ (.A(_01314_),
    .B(net271),
    .C(_01313_),
    .Y(_01316_));
 sky130_fd_sc_hd__nand3_1 _25541_ (.A(_01312_),
    .B(net271),
    .C(_01311_),
    .Y(_01317_));
 sky130_fd_sc_hd__a31o_1 _25542_ (.A1(_01314_),
    .A2(net271),
    .A3(_01313_),
    .B1(_01296_),
    .X(_01318_));
 sky130_fd_sc_hd__o221a_2 _25543_ (.A1(_05478_),
    .A2(_05479_),
    .B1(_01294_),
    .B2(net271),
    .C1(_01317_),
    .X(_01319_));
 sky130_fd_sc_hd__a211o_1 _25544_ (.A1(_01295_),
    .A2(_01316_),
    .B1(net270),
    .C1(net268),
    .X(_01320_));
 sky130_fd_sc_hd__a31o_1 _25545_ (.A1(_01314_),
    .A2(net271),
    .A3(_01313_),
    .B1(net171),
    .X(_01321_));
 sky130_fd_sc_hd__a311oi_2 _25546_ (.A1(_01314_),
    .A2(net271),
    .A3(_01313_),
    .B1(net171),
    .C1(_01296_),
    .Y(_01322_));
 sky130_fd_sc_hd__nand3_4 _25547_ (.A(_01316_),
    .B(net172),
    .C(_01295_),
    .Y(_01323_));
 sky130_fd_sc_hd__o211ai_4 _25548_ (.A1(_01294_),
    .A2(net271),
    .B1(net171),
    .C1(_01317_),
    .Y(_01324_));
 sky130_fd_sc_hd__a21oi_1 _25549_ (.A1(_00605_),
    .A2(_00976_),
    .B1(_00980_),
    .Y(_01325_));
 sky130_fd_sc_hd__a31o_1 _25550_ (.A1(_00605_),
    .A2(_00976_),
    .A3(_00979_),
    .B1(_00980_),
    .X(_01327_));
 sky130_fd_sc_hd__a31oi_2 _25551_ (.A1(_00605_),
    .A2(_00976_),
    .A3(_00979_),
    .B1(_00980_),
    .Y(_01328_));
 sky130_fd_sc_hd__a21oi_1 _25552_ (.A1(_01323_),
    .A2(_01324_),
    .B1(_01327_),
    .Y(_01329_));
 sky130_fd_sc_hd__o2bb2ai_4 _25553_ (.A1_N(_01323_),
    .A2_N(_01324_),
    .B1(_01325_),
    .B2(_00978_),
    .Y(_01330_));
 sky130_fd_sc_hd__o211a_1 _25554_ (.A1(_01296_),
    .A2(_01321_),
    .B1(_01324_),
    .C1(_01327_),
    .X(_01331_));
 sky130_fd_sc_hd__nand3_4 _25555_ (.A(_01323_),
    .B(_01324_),
    .C(_01327_),
    .Y(_01332_));
 sky130_fd_sc_hd__nand3_1 _25556_ (.A(_01330_),
    .B(_01332_),
    .C(net244),
    .Y(_01333_));
 sky130_fd_sc_hd__o22ai_1 _25557_ (.A1(net270),
    .A2(net268),
    .B1(_01329_),
    .B2(_01331_),
    .Y(_01334_));
 sky130_fd_sc_hd__a31oi_4 _25558_ (.A1(_01330_),
    .A2(_01332_),
    .A3(net244),
    .B1(_01319_),
    .Y(_01335_));
 sky130_fd_sc_hd__a31o_1 _25559_ (.A1(_01330_),
    .A2(_01332_),
    .A3(net244),
    .B1(_01319_),
    .X(_01336_));
 sky130_fd_sc_hd__o221ai_4 _25560_ (.A1(net200),
    .A2(_00618_),
    .B1(_00998_),
    .B2(_00631_),
    .C1(_00994_),
    .Y(_01338_));
 sky130_fd_sc_hd__o21ai_1 _25561_ (.A1(net175),
    .A2(_00991_),
    .B1(_01000_),
    .Y(_01339_));
 sky130_fd_sc_hd__a311oi_4 _25562_ (.A1(_01330_),
    .A2(_01332_),
    .A3(net244),
    .B1(net173),
    .C1(_01319_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand3_1 _25563_ (.A(_01333_),
    .B(net174),
    .C(_01320_),
    .Y(_01341_));
 sky130_fd_sc_hd__a2bb2oi_2 _25564_ (.A1_N(_09134_),
    .A2_N(net192),
    .B1(_01320_),
    .B2(_01333_),
    .Y(_01342_));
 sky130_fd_sc_hd__o221ai_1 _25565_ (.A1(_09134_),
    .A2(net192),
    .B1(_01318_),
    .B2(net244),
    .C1(_01334_),
    .Y(_01343_));
 sky130_fd_sc_hd__nor2_1 _25566_ (.A(_01340_),
    .B(_01342_),
    .Y(_01344_));
 sky130_fd_sc_hd__o2111ai_1 _25567_ (.A1(net177),
    .A2(_00992_),
    .B1(_01339_),
    .C1(_01341_),
    .D1(_01343_),
    .Y(_01345_));
 sky130_fd_sc_hd__o2bb2ai_1 _25568_ (.A1_N(_00994_),
    .A2_N(_01339_),
    .B1(_01340_),
    .B2(_01342_),
    .Y(_01346_));
 sky130_fd_sc_hd__o211ai_2 _25569_ (.A1(net265),
    .A2(net264),
    .B1(_01345_),
    .C1(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__o221ai_4 _25570_ (.A1(_00991_),
    .A2(net175),
    .B1(net174),
    .B2(_01335_),
    .C1(_01338_),
    .Y(_01349_));
 sky130_fd_sc_hd__o2bb2ai_1 _25571_ (.A1_N(_00995_),
    .A2_N(_01338_),
    .B1(_01340_),
    .B2(_01342_),
    .Y(_01350_));
 sky130_fd_sc_hd__o221ai_4 _25572_ (.A1(net265),
    .A2(net264),
    .B1(_01340_),
    .B2(_01349_),
    .C1(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__o21ai_4 _25573_ (.A1(net243),
    .A2(_01335_),
    .B1(_01351_),
    .Y(_01352_));
 sky130_fd_sc_hd__o31a_4 _25574_ (.A1(net265),
    .A2(net264),
    .A3(_01335_),
    .B1(_01351_),
    .X(_01353_));
 sky130_fd_sc_hd__o211ai_4 _25575_ (.A1(_01336_),
    .A2(net243),
    .B1(net175),
    .C1(_01347_),
    .Y(_01354_));
 sky130_fd_sc_hd__o211ai_4 _25576_ (.A1(net243),
    .A2(_01335_),
    .B1(net177),
    .C1(_01351_),
    .Y(_01355_));
 sky130_fd_sc_hd__nand2_2 _25577_ (.A(_01354_),
    .B(_01355_),
    .Y(_01356_));
 sky130_fd_sc_hd__o21ai_2 _25578_ (.A1(_08314_),
    .A2(_01010_),
    .B1(_01026_),
    .Y(_01357_));
 sky130_fd_sc_hd__o22ai_4 _25579_ (.A1(net200),
    .A2(_01011_),
    .B1(_01357_),
    .B2(_01023_),
    .Y(_01358_));
 sky130_fd_sc_hd__a31oi_2 _25580_ (.A1(_01015_),
    .A2(_01024_),
    .A3(_01026_),
    .B1(_01012_),
    .Y(_01360_));
 sky130_fd_sc_hd__nand3_1 _25581_ (.A(_01358_),
    .B(_01355_),
    .C(_01354_),
    .Y(_01361_));
 sky130_fd_sc_hd__a21oi_4 _25582_ (.A1(_01354_),
    .A2(_01355_),
    .B1(_01358_),
    .Y(_01362_));
 sky130_fd_sc_hd__o221ai_4 _25583_ (.A1(net200),
    .A2(_01011_),
    .B1(_01017_),
    .B2(_01029_),
    .C1(_01356_),
    .Y(_01363_));
 sky130_fd_sc_hd__o22ai_4 _25584_ (.A1(net260),
    .A2(net255),
    .B1(_01356_),
    .B2(_01360_),
    .Y(_01364_));
 sky130_fd_sc_hd__nand3_2 _25585_ (.A(net240),
    .B(_01361_),
    .C(_01363_),
    .Y(_01365_));
 sky130_fd_sc_hd__and3_1 _25586_ (.A(_01352_),
    .B(_05993_),
    .C(_05991_),
    .X(_01366_));
 sky130_fd_sc_hd__or3_2 _25587_ (.A(net260),
    .B(net255),
    .C(_01353_),
    .X(_01367_));
 sky130_fd_sc_hd__o32a_2 _25588_ (.A1(net260),
    .A2(net255),
    .A3(_01353_),
    .B1(_01362_),
    .B2(_01364_),
    .X(_01368_));
 sky130_fd_sc_hd__o22ai_4 _25589_ (.A1(net240),
    .A2(_01353_),
    .B1(_01362_),
    .B2(_01364_),
    .Y(_01369_));
 sky130_fd_sc_hd__a311o_1 _25590_ (.A1(net240),
    .A2(_01361_),
    .A3(_01363_),
    .B1(_01366_),
    .C1(_06293_),
    .X(_01371_));
 sky130_fd_sc_hd__a22oi_4 _25591_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_01365_),
    .B2(_01367_),
    .Y(_01372_));
 sky130_fd_sc_hd__o21ai_2 _25592_ (.A1(_08307_),
    .A2(net216),
    .B1(_01369_),
    .Y(_01373_));
 sky130_fd_sc_hd__o22a_1 _25593_ (.A1(_08311_),
    .A2(net215),
    .B1(_01362_),
    .B2(_01364_),
    .X(_01374_));
 sky130_fd_sc_hd__a31o_1 _25594_ (.A1(net240),
    .A2(_01361_),
    .A3(_01363_),
    .B1(_08314_),
    .X(_01375_));
 sky130_fd_sc_hd__o221a_1 _25595_ (.A1(net240),
    .A2(_01353_),
    .B1(_01362_),
    .B2(_01364_),
    .C1(net200),
    .X(_01376_));
 sky130_fd_sc_hd__o221ai_4 _25596_ (.A1(net240),
    .A2(_01353_),
    .B1(_01362_),
    .B2(_01364_),
    .C1(net200),
    .Y(_01377_));
 sky130_fd_sc_hd__a21oi_1 _25597_ (.A1(_01367_),
    .A2(_01374_),
    .B1(_01372_),
    .Y(_01378_));
 sky130_fd_sc_hd__and3_1 _25598_ (.A(_14380_),
    .B(_00296_),
    .C(_00297_),
    .X(_01379_));
 sky130_fd_sc_hd__o211a_1 _25599_ (.A1(_00649_),
    .A2(_00669_),
    .B1(_01379_),
    .C1(_00673_),
    .X(_01380_));
 sky130_fd_sc_hd__nand3_1 _25600_ (.A(_01038_),
    .B(_01379_),
    .C(_00674_),
    .Y(_01382_));
 sky130_fd_sc_hd__o211a_1 _25601_ (.A1(_01043_),
    .A2(_01037_),
    .B1(_01039_),
    .C1(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__o211ai_4 _25602_ (.A1(_01043_),
    .A2(_01037_),
    .B1(_01039_),
    .C1(_01382_),
    .Y(_01384_));
 sky130_fd_sc_hd__nand4_4 _25603_ (.A(_01380_),
    .B(_01039_),
    .C(_01038_),
    .D(_14387_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_2 _25604_ (.A(_01384_),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__a211oi_2 _25605_ (.A1(_01384_),
    .A2(_01385_),
    .B1(_01372_),
    .C1(_01376_),
    .Y(_01387_));
 sky130_fd_sc_hd__nand2_1 _25606_ (.A(_01386_),
    .B(_01378_),
    .Y(_01388_));
 sky130_fd_sc_hd__o22ai_2 _25607_ (.A1(net239),
    .A2(_06292_),
    .B1(_01378_),
    .B2(_01386_),
    .Y(_01389_));
 sky130_fd_sc_hd__nand4_2 _25608_ (.A(_01373_),
    .B(_01377_),
    .C(_01384_),
    .D(_01385_),
    .Y(_01390_));
 sky130_fd_sc_hd__a22o_1 _25609_ (.A1(_01373_),
    .A2(_01377_),
    .B1(_01384_),
    .B2(_01385_),
    .X(_01391_));
 sky130_fd_sc_hd__o221ai_1 _25610_ (.A1(net239),
    .A2(_06292_),
    .B1(_01378_),
    .B2(_01386_),
    .C1(_01388_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand3_2 _25611_ (.A(_01391_),
    .B(net214),
    .C(_01390_),
    .Y(_01394_));
 sky130_fd_sc_hd__a21oi_2 _25612_ (.A1(_01365_),
    .A2(_01367_),
    .B1(net214),
    .Y(_01395_));
 sky130_fd_sc_hd__inv_2 _25613_ (.A(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__o221a_2 _25614_ (.A1(net214),
    .A2(_01369_),
    .B1(_01387_),
    .B2(_01389_),
    .C1(_06613_),
    .X(_01397_));
 sky130_fd_sc_hd__a211o_1 _25615_ (.A1(_01394_),
    .A2(_01396_),
    .B1(net238),
    .C1(net236),
    .X(_01398_));
 sky130_fd_sc_hd__a311oi_4 _25616_ (.A1(_01391_),
    .A2(net214),
    .A3(_01390_),
    .B1(_01395_),
    .C1(_07936_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand3_4 _25617_ (.A(_01394_),
    .B(_01396_),
    .C(_07935_),
    .Y(_01400_));
 sky130_fd_sc_hd__o221ai_4 _25618_ (.A1(net214),
    .A2(_01369_),
    .B1(_01387_),
    .B2(_01389_),
    .C1(_07936_),
    .Y(_01401_));
 sky130_fd_sc_hd__a21oi_1 _25619_ (.A1(_00684_),
    .A2(_01049_),
    .B1(_01054_),
    .Y(_01402_));
 sky130_fd_sc_hd__a31oi_4 _25620_ (.A1(_00684_),
    .A2(_01049_),
    .A3(_01053_),
    .B1(_01054_),
    .Y(_01404_));
 sky130_fd_sc_hd__o2bb2ai_4 _25621_ (.A1_N(_01400_),
    .A2_N(_01401_),
    .B1(_01402_),
    .B2(_01051_),
    .Y(_01405_));
 sky130_fd_sc_hd__nand3b_4 _25622_ (.A_N(_01404_),
    .B(_01401_),
    .C(_01400_),
    .Y(_01406_));
 sky130_fd_sc_hd__nand3_1 _25623_ (.A(_01405_),
    .B(_01406_),
    .C(net209),
    .Y(_01407_));
 sky130_fd_sc_hd__a31oi_4 _25624_ (.A1(_01405_),
    .A2(_01406_),
    .A3(net209),
    .B1(_01397_),
    .Y(_01408_));
 sky130_fd_sc_hd__a31o_1 _25625_ (.A1(_01405_),
    .A2(_01406_),
    .A3(net209),
    .B1(_01397_),
    .X(_01409_));
 sky130_fd_sc_hd__o221ai_4 _25626_ (.A1(_06922_),
    .A2(_00694_),
    .B1(_01066_),
    .B2(_07246_),
    .C1(_00716_),
    .Y(_01410_));
 sky130_fd_sc_hd__a31o_1 _25627_ (.A1(_00698_),
    .A2(_00715_),
    .A3(_01068_),
    .B1(_01069_),
    .X(_01411_));
 sky130_fd_sc_hd__a311oi_4 _25628_ (.A1(_01405_),
    .A2(_01406_),
    .A3(net209),
    .B1(net202),
    .C1(_01397_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand3_2 _25629_ (.A(_01407_),
    .B(_07564_),
    .C(_01398_),
    .Y(_01413_));
 sky130_fd_sc_hd__a2bb2oi_2 _25630_ (.A1_N(net221),
    .A2_N(net220),
    .B1(_01398_),
    .B2(_01407_),
    .Y(_01415_));
 sky130_fd_sc_hd__a22o_1 _25631_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_01398_),
    .B2(_01407_),
    .X(_01416_));
 sky130_fd_sc_hd__nor2_1 _25632_ (.A(_01412_),
    .B(_01415_),
    .Y(_01417_));
 sky130_fd_sc_hd__o2111ai_2 _25633_ (.A1(_01069_),
    .A2(_01073_),
    .B1(_01413_),
    .C1(_01416_),
    .D1(_01068_),
    .Y(_01418_));
 sky130_fd_sc_hd__o221ai_4 _25634_ (.A1(net229),
    .A2(net228),
    .B1(_01411_),
    .B2(_01417_),
    .C1(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__o221ai_4 _25635_ (.A1(_01065_),
    .A2(net223),
    .B1(_07564_),
    .B2(_01408_),
    .C1(_01410_),
    .Y(_01420_));
 sky130_fd_sc_hd__o21ai_1 _25636_ (.A1(_01412_),
    .A2(_01415_),
    .B1(_01411_),
    .Y(_01421_));
 sky130_fd_sc_hd__o221ai_4 _25637_ (.A1(net229),
    .A2(net228),
    .B1(_01412_),
    .B2(_01420_),
    .C1(_01421_),
    .Y(_01422_));
 sky130_fd_sc_hd__o21ai_1 _25638_ (.A1(_06903_),
    .A2(_01408_),
    .B1(_01422_),
    .Y(_01423_));
 sky130_fd_sc_hd__o31a_1 _25639_ (.A1(net229),
    .A2(net228),
    .A3(_01408_),
    .B1(_01422_),
    .X(_01424_));
 sky130_fd_sc_hd__o211ai_4 _25640_ (.A1(_01409_),
    .A2(_06903_),
    .B1(net223),
    .C1(_01419_),
    .Y(_01426_));
 sky130_fd_sc_hd__o211a_1 _25641_ (.A1(net208),
    .A2(_01408_),
    .B1(_07246_),
    .C1(_01422_),
    .X(_01427_));
 sky130_fd_sc_hd__o211ai_4 _25642_ (.A1(_06903_),
    .A2(_01408_),
    .B1(_07246_),
    .C1(_01422_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_1 _25643_ (.A(_01426_),
    .B(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hd__a31oi_2 _25644_ (.A1(_01083_),
    .A2(_01088_),
    .A3(_01090_),
    .B1(_01081_),
    .Y(_01430_));
 sky130_fd_sc_hd__and3_1 _25645_ (.A(_01423_),
    .B(_07230_),
    .C(_07228_),
    .X(_01431_));
 sky130_fd_sc_hd__o211a_1 _25646_ (.A1(_06922_),
    .A2(_01079_),
    .B1(_01098_),
    .C1(_01429_),
    .X(_01432_));
 sky130_fd_sc_hd__o21ai_2 _25647_ (.A1(_01429_),
    .A2(_01430_),
    .B1(_07233_),
    .Y(_01433_));
 sky130_fd_sc_hd__o22ai_4 _25648_ (.A1(_07233_),
    .A2(_01424_),
    .B1(_01432_),
    .B2(_01433_),
    .Y(_01434_));
 sky130_fd_sc_hd__o22a_2 _25649_ (.A1(_07233_),
    .A2(_01424_),
    .B1(_01432_),
    .B2(_01433_),
    .X(_01435_));
 sky130_fd_sc_hd__o21ai_2 _25650_ (.A1(_06914_),
    .A2(net250),
    .B1(_01434_),
    .Y(_01437_));
 sky130_fd_sc_hd__a2bb2o_1 _25651_ (.A1_N(_01432_),
    .A2_N(_01433_),
    .B1(_06919_),
    .B2(_06921_),
    .X(_01438_));
 sky130_fd_sc_hd__o221ai_1 _25652_ (.A1(_07233_),
    .A2(_01424_),
    .B1(_01432_),
    .B2(_01433_),
    .C1(_06922_),
    .Y(_01439_));
 sky130_fd_sc_hd__o2111ai_2 _25653_ (.A1(_14451_),
    .A2(_14443_),
    .B1(_14450_),
    .C1(_00364_),
    .D1(_00366_),
    .Y(_01440_));
 sky130_fd_sc_hd__a211oi_2 _25654_ (.A1(_00720_),
    .A2(_00743_),
    .B1(_01440_),
    .C1(_00747_),
    .Y(_01441_));
 sky130_fd_sc_hd__o21ai_1 _25655_ (.A1(net233),
    .A2(_01101_),
    .B1(_01441_),
    .Y(_01442_));
 sky130_fd_sc_hd__o211ai_4 _25656_ (.A1(_01102_),
    .A2(net235),
    .B1(_01442_),
    .C1(_01114_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand4_4 _25657_ (.A(_01105_),
    .B(_01441_),
    .C(_01106_),
    .D(_14463_),
    .Y(_01444_));
 sky130_fd_sc_hd__nand2_1 _25658_ (.A(_01443_),
    .B(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__a22o_2 _25659_ (.A1(_01437_),
    .A2(_01439_),
    .B1(_01443_),
    .B2(_01444_),
    .X(_01446_));
 sky130_fd_sc_hd__o21a_1 _25660_ (.A1(net226),
    .A2(_01434_),
    .B1(_01444_),
    .X(_01448_));
 sky130_fd_sc_hd__o211ai_4 _25661_ (.A1(_01434_),
    .A2(net226),
    .B1(_01444_),
    .C1(_01443_),
    .Y(_01449_));
 sky130_fd_sc_hd__o2111ai_4 _25662_ (.A1(net226),
    .A2(_01434_),
    .B1(_01437_),
    .C1(_01443_),
    .D1(_01444_),
    .Y(_01450_));
 sky130_fd_sc_hd__nand3_2 _25663_ (.A(_01446_),
    .B(_01450_),
    .C(net163),
    .Y(_01451_));
 sky130_fd_sc_hd__and3_2 _25664_ (.A(_01434_),
    .B(_07547_),
    .C(_07545_),
    .X(_01452_));
 sky130_fd_sc_hd__or3_2 _25665_ (.A(_07544_),
    .B(_07546_),
    .C(_01435_),
    .X(_01453_));
 sky130_fd_sc_hd__a31oi_4 _25666_ (.A1(_01446_),
    .A2(_01450_),
    .A3(net163),
    .B1(_01452_),
    .Y(_01454_));
 sky130_fd_sc_hd__a21oi_1 _25667_ (.A1(_01451_),
    .A2(_01453_),
    .B1(net162),
    .Y(_01455_));
 sky130_fd_sc_hd__or3_1 _25668_ (.A(net183),
    .B(net182),
    .C(_01454_),
    .X(_01456_));
 sky130_fd_sc_hd__a31o_1 _25669_ (.A1(_01446_),
    .A2(_01450_),
    .A3(net163),
    .B1(net233),
    .X(_01457_));
 sky130_fd_sc_hd__a311oi_4 _25670_ (.A1(_01446_),
    .A2(_01450_),
    .A3(net163),
    .B1(_01452_),
    .C1(net233),
    .Y(_01459_));
 sky130_fd_sc_hd__a22oi_2 _25671_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_01451_),
    .B2(_01453_),
    .Y(_01460_));
 sky130_fd_sc_hd__a21o_1 _25672_ (.A1(_01451_),
    .A2(_01453_),
    .B1(net235),
    .X(_01461_));
 sky130_fd_sc_hd__o32a_1 _25673_ (.A1(net284),
    .A2(net281),
    .A3(_01120_),
    .B1(_01123_),
    .B2(_01127_),
    .X(_01462_));
 sky130_fd_sc_hd__a21oi_2 _25674_ (.A1(_01123_),
    .A2(_01126_),
    .B1(_01127_),
    .Y(_01463_));
 sky130_fd_sc_hd__o21a_1 _25675_ (.A1(_01459_),
    .A2(_01460_),
    .B1(_01463_),
    .X(_01464_));
 sky130_fd_sc_hd__o21ai_2 _25676_ (.A1(_01459_),
    .A2(_01460_),
    .B1(_01463_),
    .Y(_01465_));
 sky130_fd_sc_hd__o21ai_2 _25677_ (.A1(net235),
    .A2(_01454_),
    .B1(_01462_),
    .Y(_01466_));
 sky130_fd_sc_hd__o211ai_2 _25678_ (.A1(_01452_),
    .A2(_01457_),
    .B1(_01462_),
    .C1(_01461_),
    .Y(_01467_));
 sky130_fd_sc_hd__o22ai_4 _25679_ (.A1(net183),
    .A2(net182),
    .B1(_01459_),
    .B2(_01466_),
    .Y(_01468_));
 sky130_fd_sc_hd__o211ai_2 _25680_ (.A1(_01459_),
    .A2(_01466_),
    .B1(net162),
    .C1(_01465_),
    .Y(_01470_));
 sky130_fd_sc_hd__o22ai_4 _25681_ (.A1(net162),
    .A2(_01454_),
    .B1(_01464_),
    .B2(_01468_),
    .Y(_01471_));
 sky130_fd_sc_hd__and3_1 _25682_ (.A(_00775_),
    .B(_00797_),
    .C(_01141_),
    .X(_01472_));
 sky130_fd_sc_hd__o31a_1 _25683_ (.A1(_06009_),
    .A2(net287),
    .A3(_01137_),
    .B1(_01145_),
    .X(_01473_));
 sky130_fd_sc_hd__o32a_1 _25684_ (.A1(_06009_),
    .A2(net287),
    .A3(_01137_),
    .B1(_01139_),
    .B2(_01145_),
    .X(_01474_));
 sky130_fd_sc_hd__a311oi_4 _25685_ (.A1(_01465_),
    .A2(_01467_),
    .A3(net162),
    .B1(_01455_),
    .C1(net252),
    .Y(_01475_));
 sky130_fd_sc_hd__o221ai_4 _25686_ (.A1(net162),
    .A2(_01454_),
    .B1(_01464_),
    .B2(_01468_),
    .C1(_06314_),
    .Y(_01476_));
 sky130_fd_sc_hd__a22oi_4 _25687_ (.A1(_06306_),
    .A2(_06308_),
    .B1(_01456_),
    .B2(_01470_),
    .Y(_01477_));
 sky130_fd_sc_hd__o21ai_2 _25688_ (.A1(net284),
    .A2(net281),
    .B1(_01471_),
    .Y(_01478_));
 sky130_fd_sc_hd__o211ai_2 _25689_ (.A1(_01142_),
    .A2(_01472_),
    .B1(_01476_),
    .C1(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__o22ai_2 _25690_ (.A1(_01139_),
    .A2(_01473_),
    .B1(_01475_),
    .B2(_01477_),
    .Y(_01481_));
 sky130_fd_sc_hd__o211ai_4 _25691_ (.A1(_08296_),
    .A2(net179),
    .B1(_01479_),
    .C1(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__a211o_1 _25692_ (.A1(_01456_),
    .A2(_01470_),
    .B1(_08296_),
    .C1(net179),
    .X(_01483_));
 sky130_fd_sc_hd__o211ai_1 _25693_ (.A1(_01139_),
    .A2(_01473_),
    .B1(_01476_),
    .C1(_01478_),
    .Y(_01484_));
 sky130_fd_sc_hd__o22ai_1 _25694_ (.A1(_01142_),
    .A2(_01472_),
    .B1(_01475_),
    .B2(_01477_),
    .Y(_01485_));
 sky130_fd_sc_hd__o211ai_2 _25695_ (.A1(_08296_),
    .A2(net179),
    .B1(_01484_),
    .C1(_01485_),
    .Y(_01486_));
 sky130_fd_sc_hd__o21ai_4 _25696_ (.A1(net159),
    .A2(_01471_),
    .B1(_01482_),
    .Y(_01487_));
 sky130_fd_sc_hd__o211a_1 _25697_ (.A1(_01471_),
    .A2(net159),
    .B1(_06014_),
    .C1(_01482_),
    .X(_01488_));
 sky130_fd_sc_hd__o211ai_2 _25698_ (.A1(_01471_),
    .A2(net159),
    .B1(_06014_),
    .C1(_01482_),
    .Y(_01489_));
 sky130_fd_sc_hd__o211ai_4 _25699_ (.A1(net285),
    .A2(_06012_),
    .B1(_01483_),
    .C1(_01486_),
    .Y(_01490_));
 sky130_fd_sc_hd__inv_2 _25700_ (.A(_01490_),
    .Y(_01492_));
 sky130_fd_sc_hd__o31a_1 _25701_ (.A1(_05765_),
    .A2(net288),
    .A3(_01156_),
    .B1(_01164_),
    .X(_01493_));
 sky130_fd_sc_hd__a31o_1 _25702_ (.A1(_00807_),
    .A2(_01161_),
    .A3(_01163_),
    .B1(_01158_),
    .X(_01494_));
 sky130_fd_sc_hd__a22o_1 _25703_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_01483_),
    .B2(_01486_),
    .X(_01495_));
 sky130_fd_sc_hd__o2bb2ai_1 _25704_ (.A1_N(_01489_),
    .A2_N(_01490_),
    .B1(_01493_),
    .B2(_01160_),
    .Y(_01496_));
 sky130_fd_sc_hd__nand3_1 _25705_ (.A(_01489_),
    .B(_01490_),
    .C(_01494_),
    .Y(_01497_));
 sky130_fd_sc_hd__nand3_4 _25706_ (.A(_01496_),
    .B(_01497_),
    .C(net149),
    .Y(_01498_));
 sky130_fd_sc_hd__o31a_2 _25707_ (.A1(_08709_),
    .A2(_08712_),
    .A3(_01487_),
    .B1(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__a2bb2oi_4 _25708_ (.A1_N(_05760_),
    .A2_N(_05762_),
    .B1(_01495_),
    .B2(_01498_),
    .Y(_01500_));
 sky130_fd_sc_hd__o221a_1 _25709_ (.A1(_05765_),
    .A2(net288),
    .B1(net149),
    .B2(_01487_),
    .C1(_01498_),
    .X(_01501_));
 sky130_fd_sc_hd__o221ai_4 _25710_ (.A1(_05765_),
    .A2(net288),
    .B1(net149),
    .B2(_01487_),
    .C1(_01498_),
    .Y(_01503_));
 sky130_fd_sc_hd__and4_1 _25711_ (.A(_00062_),
    .B(_00064_),
    .C(_00429_),
    .D(_00431_),
    .X(_01504_));
 sky130_fd_sc_hd__nand3_1 _25712_ (.A(_00827_),
    .B(_00829_),
    .C(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__nand4_1 _25713_ (.A(_01504_),
    .B(_01179_),
    .C(_00829_),
    .D(_00827_),
    .Y(_01506_));
 sky130_fd_sc_hd__o211ai_4 _25714_ (.A1(_01177_),
    .A2(_01178_),
    .B1(_01181_),
    .C1(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hd__nand4b_2 _25715_ (.A_N(_01505_),
    .B(_01181_),
    .C(_01179_),
    .D(_00073_),
    .Y(_01508_));
 sky130_fd_sc_hd__o41ai_1 _25716_ (.A1(_00072_),
    .A2(_01178_),
    .A3(_01180_),
    .A4(_01505_),
    .B1(_01507_),
    .Y(_01509_));
 sky130_fd_sc_hd__o21ai_2 _25717_ (.A1(_01500_),
    .A2(_01501_),
    .B1(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__nand3_2 _25718_ (.A(_01503_),
    .B(_01507_),
    .C(_01508_),
    .Y(_01511_));
 sky130_fd_sc_hd__nand4b_2 _25719_ (.A_N(_01500_),
    .B(_01503_),
    .C(_01507_),
    .D(_01508_),
    .Y(_01512_));
 sky130_fd_sc_hd__o221ai_4 _25720_ (.A1(_09120_),
    .A2(net147),
    .B1(_01500_),
    .B2(_01511_),
    .C1(_01510_),
    .Y(_01514_));
 sky130_fd_sc_hd__a211o_4 _25721_ (.A1(_01495_),
    .A2(_01498_),
    .B1(net148),
    .C1(net147),
    .X(_01515_));
 sky130_fd_sc_hd__inv_2 _25722_ (.A(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__a31oi_4 _25723_ (.A1(net146),
    .A2(_01510_),
    .A3(_01512_),
    .B1(_01516_),
    .Y(_01517_));
 sky130_fd_sc_hd__a21oi_2 _25724_ (.A1(_01514_),
    .A2(_01515_),
    .B1(net143),
    .Y(_01518_));
 sky130_fd_sc_hd__or3_2 _25725_ (.A(_09553_),
    .B(net155),
    .C(_01517_),
    .X(_01519_));
 sky130_fd_sc_hd__o311a_2 _25726_ (.A1(_09120_),
    .A2(net147),
    .A3(_01499_),
    .B1(_05507_),
    .C1(_01514_),
    .X(_01520_));
 sky130_fd_sc_hd__o211ai_4 _25727_ (.A1(net146),
    .A2(_01499_),
    .B1(_05507_),
    .C1(_01514_),
    .Y(_01521_));
 sky130_fd_sc_hd__a22oi_4 _25728_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_01514_),
    .B2(_01515_),
    .Y(_01522_));
 sky130_fd_sc_hd__a22o_1 _25729_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_01514_),
    .B2(_01515_),
    .X(_01523_));
 sky130_fd_sc_hd__o21ai_2 _25730_ (.A1(_01194_),
    .A2(_01197_),
    .B1(_01193_),
    .Y(_01525_));
 sky130_fd_sc_hd__o21a_1 _25731_ (.A1(_01194_),
    .A2(_01197_),
    .B1(_01193_),
    .X(_01526_));
 sky130_fd_sc_hd__o21ai_2 _25732_ (.A1(_01520_),
    .A2(_01522_),
    .B1(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__nand3_2 _25733_ (.A(_01521_),
    .B(_01523_),
    .C(_01525_),
    .Y(_01528_));
 sky130_fd_sc_hd__o311a_1 _25734_ (.A1(_01520_),
    .A2(_01526_),
    .A3(_01522_),
    .B1(net143),
    .C1(_01527_),
    .X(_01529_));
 sky130_fd_sc_hd__nand3_4 _25735_ (.A(net143),
    .B(_01527_),
    .C(_01528_),
    .Y(_01530_));
 sky130_fd_sc_hd__o31a_1 _25736_ (.A1(_09553_),
    .A2(net155),
    .A3(_01517_),
    .B1(_01530_),
    .X(_01531_));
 sky130_fd_sc_hd__or4_1 _25737_ (.A(_09571_),
    .B(_09573_),
    .C(_01518_),
    .D(_01529_),
    .X(_01532_));
 sky130_fd_sc_hd__o21ai_2 _25738_ (.A1(_01203_),
    .A2(_01207_),
    .B1(_01202_),
    .Y(_01533_));
 sky130_fd_sc_hd__a31oi_2 _25739_ (.A1(net143),
    .A2(_01527_),
    .A3(_01528_),
    .B1(_05249_),
    .Y(_01534_));
 sky130_fd_sc_hd__o211a_1 _25740_ (.A1(net143),
    .A2(_01517_),
    .B1(_05248_),
    .C1(_01530_),
    .X(_01536_));
 sky130_fd_sc_hd__o211ai_4 _25741_ (.A1(net143),
    .A2(_01517_),
    .B1(_05248_),
    .C1(_01530_),
    .Y(_01537_));
 sky130_fd_sc_hd__a2bb2oi_4 _25742_ (.A1_N(net318),
    .A2_N(net315),
    .B1(_01519_),
    .B2(_01530_),
    .Y(_01538_));
 sky130_fd_sc_hd__o22ai_2 _25743_ (.A1(net318),
    .A2(net315),
    .B1(_01518_),
    .B2(_01529_),
    .Y(_01539_));
 sky130_fd_sc_hd__a21oi_1 _25744_ (.A1(_01519_),
    .A2(_01534_),
    .B1(_01538_),
    .Y(_01540_));
 sky130_fd_sc_hd__o2111ai_1 _25745_ (.A1(_01203_),
    .A2(_01207_),
    .B1(_01537_),
    .C1(_01539_),
    .D1(_01202_),
    .Y(_01541_));
 sky130_fd_sc_hd__o21ai_1 _25746_ (.A1(_01536_),
    .A2(_01538_),
    .B1(_01533_),
    .Y(_01542_));
 sky130_fd_sc_hd__o211ai_2 _25747_ (.A1(_09571_),
    .A2(_09573_),
    .B1(_01541_),
    .C1(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__o211a_1 _25748_ (.A1(_01518_),
    .A2(_01529_),
    .B1(_09572_),
    .C1(_09574_),
    .X(_01544_));
 sky130_fd_sc_hd__nand3_1 _25749_ (.A(_01539_),
    .B(_01533_),
    .C(_01537_),
    .Y(_01545_));
 sky130_fd_sc_hd__o21bai_2 _25750_ (.A1(_01536_),
    .A2(_01538_),
    .B1_N(_01533_),
    .Y(_01547_));
 sky130_fd_sc_hd__o211ai_2 _25751_ (.A1(_09571_),
    .A2(_09573_),
    .B1(_01545_),
    .C1(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__a31o_2 _25752_ (.A1(_09579_),
    .A2(_01545_),
    .A3(_01547_),
    .B1(_01544_),
    .X(_01549_));
 sky130_fd_sc_hd__o211ai_4 _25753_ (.A1(net340),
    .A2(_04184_),
    .B1(_01532_),
    .C1(_01543_),
    .Y(_01550_));
 sky130_fd_sc_hd__a31o_1 _25754_ (.A1(_09579_),
    .A2(_01545_),
    .A3(_01547_),
    .B1(_04238_),
    .X(_01551_));
 sky130_fd_sc_hd__o211a_1 _25755_ (.A1(_09579_),
    .A2(_01531_),
    .B1(_04227_),
    .C1(_01548_),
    .X(_01552_));
 sky130_fd_sc_hd__o211ai_4 _25756_ (.A1(_09579_),
    .A2(_01531_),
    .B1(_04227_),
    .C1(_01548_),
    .Y(_01553_));
 sky130_fd_sc_hd__a21oi_1 _25757_ (.A1(_01223_),
    .A2(_01225_),
    .B1(_01213_),
    .Y(_01554_));
 sky130_fd_sc_hd__a31oi_1 _25758_ (.A1(_01218_),
    .A2(_01223_),
    .A3(_01225_),
    .B1(_01213_),
    .Y(_01555_));
 sky130_fd_sc_hd__o2111ai_4 _25759_ (.A1(_01226_),
    .A2(_01216_),
    .B1(_01214_),
    .C1(_01553_),
    .D1(_01550_),
    .Y(_01556_));
 sky130_fd_sc_hd__a22o_1 _25760_ (.A1(_01214_),
    .A2(_01234_),
    .B1(_01550_),
    .B2(_01553_),
    .X(_01558_));
 sky130_fd_sc_hd__o211ai_4 _25761_ (.A1(_10474_),
    .A2(_10475_),
    .B1(_01556_),
    .C1(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__o311a_1 _25762_ (.A1(_09579_),
    .A2(_01518_),
    .A3(_01529_),
    .B1(_10479_),
    .C1(_01543_),
    .X(_01560_));
 sky130_fd_sc_hd__o2bb2ai_1 _25763_ (.A1_N(_01550_),
    .A2_N(_01553_),
    .B1(_01554_),
    .B2(_01216_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand3b_1 _25764_ (.A_N(_01555_),
    .B(_01553_),
    .C(_01550_),
    .Y(_01562_));
 sky130_fd_sc_hd__o211ai_1 _25765_ (.A1(_10474_),
    .A2(_10475_),
    .B1(_01561_),
    .C1(_01562_),
    .Y(_01563_));
 sky130_fd_sc_hd__o21ai_4 _25766_ (.A1(net131),
    .A2(_01549_),
    .B1(_01559_),
    .Y(_01564_));
 sky130_fd_sc_hd__o211a_1 _25767_ (.A1(_01549_),
    .A2(net131),
    .B1(_02148_),
    .C1(_01559_),
    .X(_01565_));
 sky130_fd_sc_hd__o2111ai_4 _25768_ (.A1(_01549_),
    .A2(net131),
    .B1(_02126_),
    .C1(_02104_),
    .D1(_01559_),
    .Y(_01566_));
 sky130_fd_sc_hd__nand3b_2 _25769_ (.A_N(_01560_),
    .B(_01563_),
    .C(_02137_),
    .Y(_01567_));
 sky130_fd_sc_hd__nand2_1 _25770_ (.A(_01566_),
    .B(_01567_),
    .Y(_01569_));
 sky130_fd_sc_hd__and4_1 _25771_ (.A(_00121_),
    .B(_00123_),
    .C(_00496_),
    .D(_00498_),
    .X(_01570_));
 sky130_fd_sc_hd__nand3_1 _25772_ (.A(_01240_),
    .B(_01570_),
    .C(_00887_),
    .Y(_01571_));
 sky130_fd_sc_hd__o211ai_4 _25773_ (.A1(_01237_),
    .A2(_01238_),
    .B1(_01242_),
    .C1(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand4b_1 _25774_ (.A_N(_00884_),
    .B(_01570_),
    .C(_00886_),
    .D(_00124_),
    .Y(_01573_));
 sky130_fd_sc_hd__nand3b_2 _25775_ (.A_N(_01573_),
    .B(_01242_),
    .C(_01240_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2_1 _25776_ (.A(_01572_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__or3_1 _25777_ (.A(_10949_),
    .B(net136),
    .C(_01564_),
    .X(_01576_));
 sky130_fd_sc_hd__a22o_1 _25778_ (.A1(_01566_),
    .A2(_01567_),
    .B1(_01572_),
    .B2(_01574_),
    .X(_01577_));
 sky130_fd_sc_hd__nand3_2 _25779_ (.A(_01567_),
    .B(_01572_),
    .C(_01574_),
    .Y(_01578_));
 sky130_fd_sc_hd__o221ai_4 _25780_ (.A1(_10949_),
    .A2(net136),
    .B1(_01565_),
    .B2(_01578_),
    .C1(_01577_),
    .Y(_01580_));
 sky130_fd_sc_hd__o31a_1 _25781_ (.A1(_10949_),
    .A2(net136),
    .A3(_01564_),
    .B1(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__o311a_1 _25782_ (.A1(_10949_),
    .A2(net136),
    .A3(_01564_),
    .B1(_00240_),
    .C1(_01580_),
    .X(_01582_));
 sky130_fd_sc_hd__o211ai_4 _25783_ (.A1(_10954_),
    .A2(_01564_),
    .B1(_00240_),
    .C1(_01580_),
    .Y(_01583_));
 sky130_fd_sc_hd__a22o_2 _25784_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_01576_),
    .B2(_01580_),
    .X(_01584_));
 sky130_fd_sc_hd__o32a_1 _25785_ (.A1(net361),
    .A2(net345),
    .A3(_01247_),
    .B1(_01249_),
    .B2(_01254_),
    .X(_01585_));
 sky130_fd_sc_hd__a21oi_1 _25786_ (.A1(_01254_),
    .A2(_01253_),
    .B1(_01249_),
    .Y(_01586_));
 sky130_fd_sc_hd__a21oi_1 _25787_ (.A1(_01583_),
    .A2(_01584_),
    .B1(_01585_),
    .Y(_01587_));
 sky130_fd_sc_hd__a31o_1 _25788_ (.A1(_01583_),
    .A2(_01584_),
    .A3(_01585_),
    .B1(_11464_),
    .X(_01588_));
 sky130_fd_sc_hd__o22ai_4 _25789_ (.A1(_11465_),
    .A2(_01581_),
    .B1(_01587_),
    .B2(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__o21a_1 _25790_ (.A1(net361),
    .A2(net345),
    .B1(_01589_),
    .X(_01591_));
 sky130_fd_sc_hd__o21ai_1 _25791_ (.A1(net361),
    .A2(net345),
    .B1(_01589_),
    .Y(_01592_));
 sky130_fd_sc_hd__or3_1 _25792_ (.A(net361),
    .B(net345),
    .C(_01589_),
    .X(_01593_));
 sky130_fd_sc_hd__o21ai_2 _25793_ (.A1(_01260_),
    .A2(_01262_),
    .B1(_01259_),
    .Y(_01594_));
 sky130_fd_sc_hd__a21o_1 _25794_ (.A1(_01592_),
    .A2(_01593_),
    .B1(_01594_),
    .X(_01595_));
 sky130_fd_sc_hd__a21oi_1 _25795_ (.A1(_01595_),
    .A2(_11943_),
    .B1(_01589_),
    .Y(_01596_));
 sky130_fd_sc_hd__xnor2_1 _25796_ (.A(_01265_),
    .B(_01596_),
    .Y(net100));
 sky130_fd_sc_hd__or4b_2 _25797_ (.A(_00521_),
    .B(_00908_),
    .C(_01264_),
    .D_N(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__a31o_1 _25798_ (.A1(_01567_),
    .A2(_01572_),
    .A3(_01574_),
    .B1(_01565_),
    .X(_01598_));
 sky130_fd_sc_hd__o211ai_2 _25799_ (.A1(_01266_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_01273_),
    .Y(_01599_));
 sky130_fd_sc_hd__o21ai_2 _25800_ (.A1(net304),
    .A2(_01951_),
    .B1(_01599_),
    .Y(_01601_));
 sky130_fd_sc_hd__or3_1 _25801_ (.A(net302),
    .B(_04019_),
    .C(_01601_),
    .X(_01602_));
 sky130_fd_sc_hd__a21o_1 _25802_ (.A1(_10963_),
    .A2(_10964_),
    .B1(_01601_),
    .X(_01603_));
 sky130_fd_sc_hd__a22o_1 _25803_ (.A1(_10966_),
    .A2(_10968_),
    .B1(_01599_),
    .B2(net278),
    .X(_01604_));
 sky130_fd_sc_hd__xor2_1 _25804_ (.A(_10970_),
    .B(_01601_),
    .X(_01605_));
 sky130_fd_sc_hd__nand2_1 _25805_ (.A(_01603_),
    .B(_01604_),
    .Y(_01606_));
 sky130_fd_sc_hd__o21ai_1 _25806_ (.A1(_01281_),
    .A2(_01286_),
    .B1(_01279_),
    .Y(_01607_));
 sky130_fd_sc_hd__nand2_1 _25807_ (.A(_01607_),
    .B(_01605_),
    .Y(_01608_));
 sky130_fd_sc_hd__o211ai_1 _25808_ (.A1(_01286_),
    .A2(_01285_),
    .B1(_01279_),
    .C1(_01606_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand3_2 _25809_ (.A(_01608_),
    .B(_01609_),
    .C(_04029_),
    .Y(_01610_));
 sky130_fd_sc_hd__a21oi_1 _25810_ (.A1(_01602_),
    .A2(_01610_),
    .B1(net150),
    .Y(_01612_));
 sky130_fd_sc_hd__a2bb2o_2 _25811_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_01602_),
    .B2(_01610_),
    .X(_01613_));
 sky130_fd_sc_hd__and3_1 _25812_ (.A(_01610_),
    .B(net150),
    .C(_01602_),
    .X(_01614_));
 sky130_fd_sc_hd__o211ai_2 _25813_ (.A1(_04029_),
    .A2(_01601_),
    .B1(net150),
    .C1(_01610_),
    .Y(_01615_));
 sky130_fd_sc_hd__a22o_1 _25814_ (.A1(net151),
    .A2(_01294_),
    .B1(_01308_),
    .B2(_01309_),
    .X(_01616_));
 sky130_fd_sc_hd__a31oi_2 _25815_ (.A1(_01300_),
    .A2(_01308_),
    .A3(_01309_),
    .B1(_01297_),
    .Y(_01617_));
 sky130_fd_sc_hd__o21ai_2 _25816_ (.A1(_01612_),
    .A2(_01614_),
    .B1(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__o2111ai_4 _25817_ (.A1(net151),
    .A2(_01294_),
    .B1(_01613_),
    .C1(_01615_),
    .D1(_01616_),
    .Y(_01619_));
 sky130_fd_sc_hd__a211o_2 _25818_ (.A1(_01602_),
    .A2(_01610_),
    .B1(net296),
    .C1(_05232_),
    .X(_01620_));
 sky130_fd_sc_hd__inv_2 _25819_ (.A(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__o211a_1 _25820_ (.A1(net296),
    .A2(_05232_),
    .B1(_01618_),
    .C1(_01619_),
    .X(_01623_));
 sky130_fd_sc_hd__o211ai_4 _25821_ (.A1(net296),
    .A2(_05232_),
    .B1(_01618_),
    .C1(_01619_),
    .Y(_01624_));
 sky130_fd_sc_hd__nor2_1 _25822_ (.A(_01621_),
    .B(_01623_),
    .Y(_01625_));
 sky130_fd_sc_hd__o22a_2 _25823_ (.A1(_05478_),
    .A2(_05479_),
    .B1(_01621_),
    .B2(_01623_),
    .X(_01626_));
 sky130_fd_sc_hd__a211o_1 _25824_ (.A1(_01620_),
    .A2(_01624_),
    .B1(net270),
    .C1(net268),
    .X(_01627_));
 sky130_fd_sc_hd__and3_1 _25825_ (.A(_00245_),
    .B(_00603_),
    .C(_00605_),
    .X(_01628_));
 sky130_fd_sc_hd__nand3_1 _25826_ (.A(_01323_),
    .B(_01628_),
    .C(_00982_),
    .Y(_01629_));
 sky130_fd_sc_hd__o211ai_4 _25827_ (.A1(_01328_),
    .A2(_01322_),
    .B1(_01324_),
    .C1(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__nand4_1 _25828_ (.A(_01628_),
    .B(_00981_),
    .C(_00979_),
    .D(_00254_),
    .Y(_01631_));
 sky130_fd_sc_hd__nand4_4 _25829_ (.A(_01323_),
    .B(_01324_),
    .C(_01628_),
    .D(_00982_),
    .Y(_01632_));
 sky130_fd_sc_hd__nand3b_4 _25830_ (.A_N(_01631_),
    .B(_01324_),
    .C(_01323_),
    .Y(_01634_));
 sky130_fd_sc_hd__o21ai_1 _25831_ (.A1(_00255_),
    .A2(_01632_),
    .B1(_01630_),
    .Y(_01635_));
 sky130_fd_sc_hd__a31oi_1 _25832_ (.A1(_01618_),
    .A2(_01619_),
    .A3(net271),
    .B1(net151),
    .Y(_01636_));
 sky130_fd_sc_hd__and3_1 _25833_ (.A(_01624_),
    .B(net153),
    .C(_01620_),
    .X(_01637_));
 sky130_fd_sc_hd__o211ai_4 _25834_ (.A1(net167),
    .A2(_10024_),
    .B1(_01620_),
    .C1(_01624_),
    .Y(_01638_));
 sky130_fd_sc_hd__a2bb2oi_4 _25835_ (.A1_N(net170),
    .A2_N(_10022_),
    .B1(_01620_),
    .B2(_01624_),
    .Y(_01639_));
 sky130_fd_sc_hd__o22ai_2 _25836_ (.A1(net170),
    .A2(_10022_),
    .B1(_01621_),
    .B2(_01623_),
    .Y(_01640_));
 sky130_fd_sc_hd__a21oi_1 _25837_ (.A1(_01620_),
    .A2(_01636_),
    .B1(_01639_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_1 _25838_ (.A(_01635_),
    .B(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__o221ai_2 _25839_ (.A1(_01632_),
    .A2(_00255_),
    .B1(_01639_),
    .B2(_01637_),
    .C1(_01630_),
    .Y(_01643_));
 sky130_fd_sc_hd__o2bb2ai_2 _25840_ (.A1_N(_01630_),
    .A2_N(_01634_),
    .B1(_01637_),
    .B2(_01639_),
    .Y(_01645_));
 sky130_fd_sc_hd__o2111ai_4 _25841_ (.A1(_00255_),
    .A2(_01632_),
    .B1(_01638_),
    .C1(_01640_),
    .D1(_01630_),
    .Y(_01646_));
 sky130_fd_sc_hd__nand3_1 _25842_ (.A(_01645_),
    .B(_01646_),
    .C(net244),
    .Y(_01647_));
 sky130_fd_sc_hd__or4_1 _25843_ (.A(net270),
    .B(net268),
    .C(_01621_),
    .D(_01623_),
    .X(_01648_));
 sky130_fd_sc_hd__nand3_2 _25844_ (.A(_01642_),
    .B(_01643_),
    .C(net244),
    .Y(_01649_));
 sky130_fd_sc_hd__a31o_1 _25845_ (.A1(_01645_),
    .A2(_01646_),
    .A3(net244),
    .B1(_01626_),
    .X(_01650_));
 sky130_fd_sc_hd__o311a_2 _25846_ (.A1(net244),
    .A2(_01621_),
    .A3(_01623_),
    .B1(_01649_),
    .C1(_05754_),
    .X(_01651_));
 sky130_fd_sc_hd__a211o_2 _25847_ (.A1(_01627_),
    .A2(_01647_),
    .B1(net265),
    .C1(net264),
    .X(_01652_));
 sky130_fd_sc_hd__a31o_1 _25848_ (.A1(_01645_),
    .A2(_01646_),
    .A3(net244),
    .B1(net171),
    .X(_01653_));
 sky130_fd_sc_hd__a311oi_2 _25849_ (.A1(_01645_),
    .A2(_01646_),
    .A3(net244),
    .B1(net171),
    .C1(_01626_),
    .Y(_01654_));
 sky130_fd_sc_hd__nand3_4 _25850_ (.A(_01647_),
    .B(net172),
    .C(_01627_),
    .Y(_01656_));
 sky130_fd_sc_hd__o211ai_4 _25851_ (.A1(net189),
    .A2(net188),
    .B1(_01648_),
    .C1(_01649_),
    .Y(_01657_));
 sky130_fd_sc_hd__o221a_1 _25852_ (.A1(net177),
    .A2(_00992_),
    .B1(_01335_),
    .B2(net174),
    .C1(_01339_),
    .X(_01658_));
 sky130_fd_sc_hd__a31o_1 _25853_ (.A1(_00995_),
    .A2(_01338_),
    .A3(_01341_),
    .B1(_01342_),
    .X(_01659_));
 sky130_fd_sc_hd__a31oi_2 _25854_ (.A1(_00995_),
    .A2(_01338_),
    .A3(_01341_),
    .B1(_01342_),
    .Y(_01660_));
 sky130_fd_sc_hd__a21oi_1 _25855_ (.A1(_01656_),
    .A2(_01657_),
    .B1(_01659_),
    .Y(_01661_));
 sky130_fd_sc_hd__o2bb2ai_4 _25856_ (.A1_N(_01656_),
    .A2_N(_01657_),
    .B1(_01658_),
    .B2(_01340_),
    .Y(_01662_));
 sky130_fd_sc_hd__o211a_1 _25857_ (.A1(_01626_),
    .A2(_01653_),
    .B1(_01657_),
    .C1(_01659_),
    .X(_01663_));
 sky130_fd_sc_hd__o211ai_4 _25858_ (.A1(_01626_),
    .A2(_01653_),
    .B1(_01657_),
    .C1(_01659_),
    .Y(_01664_));
 sky130_fd_sc_hd__nand3_2 _25859_ (.A(_01662_),
    .B(_01664_),
    .C(net243),
    .Y(_01665_));
 sky130_fd_sc_hd__o22ai_1 _25860_ (.A1(net265),
    .A2(net264),
    .B1(_01661_),
    .B2(_01663_),
    .Y(_01667_));
 sky130_fd_sc_hd__a31oi_4 _25861_ (.A1(_01662_),
    .A2(_01664_),
    .A3(net243),
    .B1(_01651_),
    .Y(_01668_));
 sky130_fd_sc_hd__a311o_1 _25862_ (.A1(_01662_),
    .A2(_01664_),
    .A3(net243),
    .B1(net240),
    .C1(_01651_),
    .X(_01669_));
 sky130_fd_sc_hd__o221ai_4 _25863_ (.A1(net200),
    .A2(_01011_),
    .B1(_01357_),
    .B2(_01023_),
    .C1(_01354_),
    .Y(_01670_));
 sky130_fd_sc_hd__o21ai_1 _25864_ (.A1(_08731_),
    .A2(_01352_),
    .B1(_01358_),
    .Y(_01671_));
 sky130_fd_sc_hd__a31oi_2 _25865_ (.A1(_01662_),
    .A2(_01664_),
    .A3(net243),
    .B1(net173),
    .Y(_01672_));
 sky130_fd_sc_hd__a311oi_4 _25866_ (.A1(_01662_),
    .A2(_01664_),
    .A3(net243),
    .B1(net173),
    .C1(_01651_),
    .Y(_01673_));
 sky130_fd_sc_hd__nand3_2 _25867_ (.A(_01665_),
    .B(net174),
    .C(_01652_),
    .Y(_01674_));
 sky130_fd_sc_hd__a2bb2oi_4 _25868_ (.A1_N(net194),
    .A2_N(net192),
    .B1(_01652_),
    .B2(_01665_),
    .Y(_01675_));
 sky130_fd_sc_hd__o221ai_1 _25869_ (.A1(net194),
    .A2(net192),
    .B1(_01650_),
    .B2(_05752_),
    .C1(_01667_),
    .Y(_01676_));
 sky130_fd_sc_hd__a21oi_1 _25870_ (.A1(_01652_),
    .A2(_01672_),
    .B1(_01675_),
    .Y(_01678_));
 sky130_fd_sc_hd__o2111ai_1 _25871_ (.A1(net177),
    .A2(_01353_),
    .B1(_01671_),
    .C1(_01674_),
    .D1(_01676_),
    .Y(_01679_));
 sky130_fd_sc_hd__o2bb2ai_1 _25872_ (.A1_N(_01354_),
    .A2_N(_01671_),
    .B1(_01673_),
    .B2(_01675_),
    .Y(_01680_));
 sky130_fd_sc_hd__nand3_1 _25873_ (.A(net240),
    .B(_01679_),
    .C(_01680_),
    .Y(_01681_));
 sky130_fd_sc_hd__or3_1 _25874_ (.A(net260),
    .B(net255),
    .C(_01668_),
    .X(_01682_));
 sky130_fd_sc_hd__o221ai_4 _25875_ (.A1(_01352_),
    .A2(_08731_),
    .B1(net174),
    .B2(_01668_),
    .C1(_01670_),
    .Y(_01683_));
 sky130_fd_sc_hd__o2bb2ai_1 _25876_ (.A1_N(_01355_),
    .A2_N(_01670_),
    .B1(_01673_),
    .B2(_01675_),
    .Y(_01684_));
 sky130_fd_sc_hd__o221ai_4 _25877_ (.A1(net260),
    .A2(net255),
    .B1(_01673_),
    .B2(_01683_),
    .C1(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__o21ai_2 _25878_ (.A1(net240),
    .A2(_01668_),
    .B1(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__o221a_2 _25879_ (.A1(_06286_),
    .A2(_06288_),
    .B1(_01668_),
    .B2(net240),
    .C1(_01685_),
    .X(_01687_));
 sky130_fd_sc_hd__a2bb2oi_2 _25880_ (.A1_N(_08724_),
    .A2_N(net196),
    .B1(_01682_),
    .B2(_01685_),
    .Y(_01689_));
 sky130_fd_sc_hd__o211ai_4 _25881_ (.A1(_08724_),
    .A2(net196),
    .B1(_01669_),
    .C1(_01681_),
    .Y(_01690_));
 sky130_fd_sc_hd__o311a_1 _25882_ (.A1(net260),
    .A2(net255),
    .A3(_01668_),
    .B1(net178),
    .C1(_01685_),
    .X(_01691_));
 sky130_fd_sc_hd__o211ai_4 _25883_ (.A1(net240),
    .A2(_01668_),
    .B1(net178),
    .C1(_01685_),
    .Y(_01692_));
 sky130_fd_sc_hd__nand2_1 _25884_ (.A(_01690_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__o21ai_2 _25885_ (.A1(_08314_),
    .A2(_01369_),
    .B1(_01385_),
    .Y(_01694_));
 sky130_fd_sc_hd__o211ai_2 _25886_ (.A1(_01375_),
    .A2(_01366_),
    .B1(_01385_),
    .C1(_01384_),
    .Y(_01695_));
 sky130_fd_sc_hd__o22ai_2 _25887_ (.A1(net200),
    .A2(_01368_),
    .B1(_01694_),
    .B2(_01383_),
    .Y(_01696_));
 sky130_fd_sc_hd__a31oi_2 _25888_ (.A1(_01377_),
    .A2(_01384_),
    .A3(_01385_),
    .B1(_01372_),
    .Y(_01697_));
 sky130_fd_sc_hd__o2111ai_4 _25889_ (.A1(net200),
    .A2(_01368_),
    .B1(_01690_),
    .C1(_01692_),
    .D1(_01695_),
    .Y(_01698_));
 sky130_fd_sc_hd__o21ai_2 _25890_ (.A1(_01689_),
    .A2(_01691_),
    .B1(_01696_),
    .Y(_01700_));
 sky130_fd_sc_hd__o211ai_1 _25891_ (.A1(net239),
    .A2(_06292_),
    .B1(_01698_),
    .C1(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__a22o_1 _25892_ (.A1(_06287_),
    .A2(_06290_),
    .B1(_01682_),
    .B2(_01685_),
    .X(_01702_));
 sky130_fd_sc_hd__nand3_1 _25893_ (.A(_01696_),
    .B(_01692_),
    .C(_01690_),
    .Y(_01703_));
 sky130_fd_sc_hd__a21oi_1 _25894_ (.A1(_01690_),
    .A2(_01692_),
    .B1(_01696_),
    .Y(_01704_));
 sky130_fd_sc_hd__o21ai_1 _25895_ (.A1(_01689_),
    .A2(_01691_),
    .B1(_01697_),
    .Y(_01705_));
 sky130_fd_sc_hd__o22ai_2 _25896_ (.A1(net239),
    .A2(_06292_),
    .B1(_01693_),
    .B2(_01697_),
    .Y(_01706_));
 sky130_fd_sc_hd__a31o_2 _25897_ (.A1(_01700_),
    .A2(net214),
    .A3(_01698_),
    .B1(_01687_),
    .X(_01707_));
 sky130_fd_sc_hd__inv_2 _25898_ (.A(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__a311oi_4 _25899_ (.A1(_01700_),
    .A2(net214),
    .A3(_01698_),
    .B1(net200),
    .C1(_01687_),
    .Y(_01709_));
 sky130_fd_sc_hd__o211ai_1 _25900_ (.A1(net214),
    .A2(_01686_),
    .B1(_01701_),
    .C1(_08314_),
    .Y(_01711_));
 sky130_fd_sc_hd__a31oi_1 _25901_ (.A1(_01703_),
    .A2(_01705_),
    .A3(_06293_),
    .B1(_08314_),
    .Y(_01712_));
 sky130_fd_sc_hd__o211ai_4 _25902_ (.A1(_01704_),
    .A2(_01706_),
    .B1(net200),
    .C1(_01702_),
    .Y(_01713_));
 sky130_fd_sc_hd__a21oi_2 _25903_ (.A1(_01712_),
    .A2(_01702_),
    .B1(_01709_),
    .Y(_01714_));
 sky130_fd_sc_hd__nand2_1 _25904_ (.A(_01711_),
    .B(_01713_),
    .Y(_01715_));
 sky130_fd_sc_hd__o2111a_1 _25905_ (.A1(_00310_),
    .A2(_00303_),
    .B1(_00309_),
    .C1(_00684_),
    .D1(_00685_),
    .X(_01716_));
 sky130_fd_sc_hd__o2111ai_1 _25906_ (.A1(_00310_),
    .A2(_00303_),
    .B1(_00309_),
    .C1(_00684_),
    .D1(_00685_),
    .Y(_01717_));
 sky130_fd_sc_hd__o21ai_1 _25907_ (.A1(_07564_),
    .A2(_01047_),
    .B1(_01716_),
    .Y(_01718_));
 sky130_fd_sc_hd__nor3_1 _25908_ (.A(_01051_),
    .B(_01717_),
    .C(_01054_),
    .Y(_01719_));
 sky130_fd_sc_hd__nand2_1 _25909_ (.A(_01400_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__a32oi_1 _25910_ (.A1(_07936_),
    .A2(_01371_),
    .A3(_01393_),
    .B1(_01400_),
    .B2(_01719_),
    .Y(_01722_));
 sky130_fd_sc_hd__o311a_1 _25911_ (.A1(_01051_),
    .A2(_01718_),
    .A3(_01399_),
    .B1(_01401_),
    .C1(_01406_),
    .X(_01723_));
 sky130_fd_sc_hd__o211ai_4 _25912_ (.A1(_01404_),
    .A2(_01399_),
    .B1(_01401_),
    .C1(_01720_),
    .Y(_01724_));
 sky130_fd_sc_hd__nor3_1 _25913_ (.A(_00318_),
    .B(_01051_),
    .C(_01718_),
    .Y(_01725_));
 sky130_fd_sc_hd__nand3_4 _25914_ (.A(_01725_),
    .B(_01401_),
    .C(_01400_),
    .Y(_01726_));
 sky130_fd_sc_hd__a21boi_1 _25915_ (.A1(_01722_),
    .A2(_01406_),
    .B1_N(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__nand2_1 _25916_ (.A(_01724_),
    .B(_01726_),
    .Y(_01728_));
 sky130_fd_sc_hd__a21oi_2 _25917_ (.A1(_01724_),
    .A2(_01726_),
    .B1(_01715_),
    .Y(_01729_));
 sky130_fd_sc_hd__a31o_1 _25918_ (.A1(_01715_),
    .A2(_01724_),
    .A3(_01726_),
    .B1(_06613_),
    .X(_01730_));
 sky130_fd_sc_hd__nand3_2 _25919_ (.A(_01714_),
    .B(_01724_),
    .C(_01726_),
    .Y(_01731_));
 sky130_fd_sc_hd__a22o_1 _25920_ (.A1(_01711_),
    .A2(_01713_),
    .B1(_01724_),
    .B2(_01726_),
    .X(_01733_));
 sky130_fd_sc_hd__o221ai_4 _25921_ (.A1(net238),
    .A2(net236),
    .B1(_01714_),
    .B2(_01727_),
    .C1(_01731_),
    .Y(_01734_));
 sky130_fd_sc_hd__o211a_1 _25922_ (.A1(net214),
    .A2(_01686_),
    .B1(_01701_),
    .C1(_06613_),
    .X(_01735_));
 sky130_fd_sc_hd__a311o_1 _25923_ (.A1(_01700_),
    .A2(net214),
    .A3(_01698_),
    .B1(net209),
    .C1(_01687_),
    .X(_01736_));
 sky130_fd_sc_hd__o221a_1 _25924_ (.A1(net209),
    .A2(_01708_),
    .B1(_01729_),
    .B2(_01730_),
    .C1(_06904_),
    .X(_01737_));
 sky130_fd_sc_hd__a211o_2 _25925_ (.A1(_01734_),
    .A2(_01736_),
    .B1(net229),
    .C1(net228),
    .X(_01738_));
 sky130_fd_sc_hd__a311oi_4 _25926_ (.A1(_01733_),
    .A2(net209),
    .A3(_01731_),
    .B1(_01735_),
    .C1(_07936_),
    .Y(_01739_));
 sky130_fd_sc_hd__nand3_4 _25927_ (.A(_01734_),
    .B(_01736_),
    .C(_07935_),
    .Y(_01740_));
 sky130_fd_sc_hd__o221ai_4 _25928_ (.A1(net209),
    .A2(_01708_),
    .B1(_01729_),
    .B2(_01730_),
    .C1(_07936_),
    .Y(_01741_));
 sky130_fd_sc_hd__o221a_1 _25929_ (.A1(_07564_),
    .A2(_01408_),
    .B1(_01073_),
    .B2(_01069_),
    .C1(_01068_),
    .X(_01742_));
 sky130_fd_sc_hd__a31o_1 _25930_ (.A1(_01070_),
    .A2(_01410_),
    .A3(_01413_),
    .B1(_01415_),
    .X(_01744_));
 sky130_fd_sc_hd__a31oi_2 _25931_ (.A1(_01070_),
    .A2(_01410_),
    .A3(_01413_),
    .B1(_01415_),
    .Y(_01745_));
 sky130_fd_sc_hd__o2bb2ai_4 _25932_ (.A1_N(_01740_),
    .A2_N(_01741_),
    .B1(_01742_),
    .B2(_01412_),
    .Y(_01746_));
 sky130_fd_sc_hd__nand3_2 _25933_ (.A(_01744_),
    .B(_01741_),
    .C(_01740_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand3_2 _25934_ (.A(_01746_),
    .B(_01747_),
    .C(_06903_),
    .Y(_01748_));
 sky130_fd_sc_hd__a31o_1 _25935_ (.A1(_01746_),
    .A2(_01747_),
    .A3(_06903_),
    .B1(_01737_),
    .X(_01749_));
 sky130_fd_sc_hd__a311o_1 _25936_ (.A1(_01746_),
    .A2(_01747_),
    .A3(_06903_),
    .B1(_07233_),
    .C1(_01737_),
    .X(_01750_));
 sky130_fd_sc_hd__a31oi_2 _25937_ (.A1(_01746_),
    .A2(_01747_),
    .A3(_06903_),
    .B1(net202),
    .Y(_01751_));
 sky130_fd_sc_hd__a311oi_2 _25938_ (.A1(_01746_),
    .A2(_01747_),
    .A3(_06903_),
    .B1(net202),
    .C1(_01737_),
    .Y(_01752_));
 sky130_fd_sc_hd__nand3_2 _25939_ (.A(_01748_),
    .B(_07564_),
    .C(_01738_),
    .Y(_01753_));
 sky130_fd_sc_hd__a2bb2oi_4 _25940_ (.A1_N(net221),
    .A2_N(net220),
    .B1(_01738_),
    .B2(_01748_),
    .Y(_01755_));
 sky130_fd_sc_hd__a22o_1 _25941_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_01738_),
    .B2(_01748_),
    .X(_01756_));
 sky130_fd_sc_hd__a21oi_1 _25942_ (.A1(_01738_),
    .A2(_01751_),
    .B1(_01755_),
    .Y(_01757_));
 sky130_fd_sc_hd__o211ai_4 _25943_ (.A1(_01079_),
    .A2(_06922_),
    .B1(_01426_),
    .C1(_01098_),
    .Y(_01758_));
 sky130_fd_sc_hd__a31o_1 _25944_ (.A1(_01082_),
    .A2(_01098_),
    .A3(_01426_),
    .B1(_01427_),
    .X(_01759_));
 sky130_fd_sc_hd__o2111ai_2 _25945_ (.A1(_01427_),
    .A2(_01430_),
    .B1(_01753_),
    .C1(_01756_),
    .D1(_01426_),
    .Y(_01760_));
 sky130_fd_sc_hd__o221ai_4 _25946_ (.A1(net207),
    .A2(net205),
    .B1(_01759_),
    .B2(_01757_),
    .C1(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__a211o_1 _25947_ (.A1(_01738_),
    .A2(_01748_),
    .B1(net207),
    .C1(net205),
    .X(_01762_));
 sky130_fd_sc_hd__o21ai_1 _25948_ (.A1(_01752_),
    .A2(_01755_),
    .B1(_01759_),
    .Y(_01763_));
 sky130_fd_sc_hd__o2111ai_1 _25949_ (.A1(net223),
    .A2(_01423_),
    .B1(_01753_),
    .C1(_01756_),
    .D1(_01758_),
    .Y(_01764_));
 sky130_fd_sc_hd__o211ai_2 _25950_ (.A1(net207),
    .A2(net205),
    .B1(_01763_),
    .C1(_01764_),
    .Y(_01766_));
 sky130_fd_sc_hd__o21ai_4 _25951_ (.A1(_07233_),
    .A2(_01749_),
    .B1(_01761_),
    .Y(_01767_));
 sky130_fd_sc_hd__o211ai_4 _25952_ (.A1(_07242_),
    .A2(net248),
    .B1(_01750_),
    .C1(_01761_),
    .Y(_01768_));
 sky130_fd_sc_hd__and3_1 _25953_ (.A(_01766_),
    .B(_07246_),
    .C(_01762_),
    .X(_01769_));
 sky130_fd_sc_hd__o211ai_4 _25954_ (.A1(_07244_),
    .A2(net247),
    .B1(_01762_),
    .C1(_01766_),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_1 _25955_ (.A(_01768_),
    .B(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__o2bb2ai_1 _25956_ (.A1_N(_01443_),
    .A2_N(_01444_),
    .B1(_06922_),
    .B2(_01435_),
    .Y(_01772_));
 sky130_fd_sc_hd__a22oi_4 _25957_ (.A1(net226),
    .A2(_01434_),
    .B1(_01448_),
    .B2(_01443_),
    .Y(_01773_));
 sky130_fd_sc_hd__o311a_1 _25958_ (.A1(_06918_),
    .A2(net249),
    .A3(_01435_),
    .B1(_01449_),
    .C1(_01771_),
    .X(_01774_));
 sky130_fd_sc_hd__o211ai_1 _25959_ (.A1(_06922_),
    .A2(_01435_),
    .B1(_01449_),
    .C1(_01771_),
    .Y(_01775_));
 sky130_fd_sc_hd__o2111ai_1 _25960_ (.A1(net226),
    .A2(_01434_),
    .B1(_01768_),
    .C1(_01770_),
    .D1(_01772_),
    .Y(_01777_));
 sky130_fd_sc_hd__o22ai_2 _25961_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_01771_),
    .B2(_01773_),
    .Y(_01778_));
 sky130_fd_sc_hd__nand3_2 _25962_ (.A(_01777_),
    .B(net163),
    .C(_01775_),
    .Y(_01779_));
 sky130_fd_sc_hd__or3_1 _25963_ (.A(_07544_),
    .B(_07546_),
    .C(_01767_),
    .X(_01780_));
 sky130_fd_sc_hd__o32a_1 _25964_ (.A1(_07544_),
    .A2(_07546_),
    .A3(_01767_),
    .B1(_01774_),
    .B2(_01778_),
    .X(_01781_));
 sky130_fd_sc_hd__o22ai_4 _25965_ (.A1(net163),
    .A2(_01767_),
    .B1(_01774_),
    .B2(_01778_),
    .Y(_01782_));
 sky130_fd_sc_hd__a22oi_2 _25966_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_01779_),
    .B2(_01780_),
    .Y(_01783_));
 sky130_fd_sc_hd__o21ai_4 _25967_ (.A1(_06914_),
    .A2(net250),
    .B1(_01782_),
    .Y(_01784_));
 sky130_fd_sc_hd__o221a_1 _25968_ (.A1(_06918_),
    .A2(net249),
    .B1(net163),
    .B2(_01767_),
    .C1(_01779_),
    .X(_01785_));
 sky130_fd_sc_hd__o221ai_4 _25969_ (.A1(_06918_),
    .A2(net249),
    .B1(net163),
    .B2(_01767_),
    .C1(_01779_),
    .Y(_01786_));
 sky130_fd_sc_hd__nand2_1 _25970_ (.A(_01784_),
    .B(_01786_),
    .Y(_01788_));
 sky130_fd_sc_hd__o2111a_1 _25971_ (.A1(_00380_),
    .A2(_00374_),
    .B1(_00379_),
    .C1(_00760_),
    .D1(_00762_),
    .X(_01789_));
 sky130_fd_sc_hd__o211ai_2 _25972_ (.A1(_01103_),
    .A2(_01124_),
    .B1(_01789_),
    .C1(_01128_),
    .Y(_01790_));
 sky130_fd_sc_hd__a31oi_2 _25973_ (.A1(_01451_),
    .A2(_01453_),
    .A3(net235),
    .B1(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__a31o_1 _25974_ (.A1(_01451_),
    .A2(_01453_),
    .A3(net235),
    .B1(_01790_),
    .X(_01792_));
 sky130_fd_sc_hd__o211ai_4 _25975_ (.A1(_01463_),
    .A2(_01459_),
    .B1(_01461_),
    .C1(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__o211ai_4 _25976_ (.A1(net235),
    .A2(_01454_),
    .B1(_00386_),
    .C1(_01791_),
    .Y(_01794_));
 sky130_fd_sc_hd__nand2_1 _25977_ (.A(_01793_),
    .B(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__a21oi_2 _25978_ (.A1(_01793_),
    .A2(_01794_),
    .B1(_01788_),
    .Y(_01796_));
 sky130_fd_sc_hd__o211ai_1 _25979_ (.A1(_01783_),
    .A2(_01785_),
    .B1(_01793_),
    .C1(_01794_),
    .Y(_01797_));
 sky130_fd_sc_hd__o21ai_2 _25980_ (.A1(net183),
    .A2(net182),
    .B1(_01797_),
    .Y(_01799_));
 sky130_fd_sc_hd__and3_1 _25981_ (.A(_07913_),
    .B(_07915_),
    .C(_01782_),
    .X(_01800_));
 sky130_fd_sc_hd__or3_2 _25982_ (.A(net183),
    .B(net182),
    .C(_01781_),
    .X(_01801_));
 sky130_fd_sc_hd__a22o_1 _25983_ (.A1(_01784_),
    .A2(_01786_),
    .B1(_01793_),
    .B2(_01794_),
    .X(_01802_));
 sky130_fd_sc_hd__nand3_2 _25984_ (.A(_01786_),
    .B(_01793_),
    .C(_01794_),
    .Y(_01803_));
 sky130_fd_sc_hd__nand4_2 _25985_ (.A(_01784_),
    .B(_01786_),
    .C(_01793_),
    .D(_01794_),
    .Y(_01804_));
 sky130_fd_sc_hd__nand3_2 _25986_ (.A(_01802_),
    .B(_01804_),
    .C(net162),
    .Y(_01805_));
 sky130_fd_sc_hd__o221a_1 _25987_ (.A1(net162),
    .A2(_01782_),
    .B1(_01796_),
    .B2(_01799_),
    .C1(_08301_),
    .X(_01806_));
 sky130_fd_sc_hd__a211o_1 _25988_ (.A1(_01801_),
    .A2(_01805_),
    .B1(_08296_),
    .C1(net179),
    .X(_01807_));
 sky130_fd_sc_hd__a311oi_4 _25989_ (.A1(_01802_),
    .A2(_01804_),
    .A3(net162),
    .B1(_01800_),
    .C1(net233),
    .Y(_01808_));
 sky130_fd_sc_hd__nand3_4 _25990_ (.A(_01805_),
    .B(net235),
    .C(_01801_),
    .Y(_01810_));
 sky130_fd_sc_hd__o221ai_4 _25991_ (.A1(net162),
    .A2(_01782_),
    .B1(_01796_),
    .B2(_01799_),
    .C1(net233),
    .Y(_01811_));
 sky130_fd_sc_hd__nand2_1 _25992_ (.A(_01810_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__o2bb2a_1 _25993_ (.A1_N(net252),
    .A2_N(_01471_),
    .B1(_01472_),
    .B2(_01142_),
    .X(_01813_));
 sky130_fd_sc_hd__a31o_1 _25994_ (.A1(_06311_),
    .A2(_06313_),
    .A3(_01471_),
    .B1(_01474_),
    .X(_01814_));
 sky130_fd_sc_hd__a21oi_2 _25995_ (.A1(_01474_),
    .A2(_01476_),
    .B1(_01477_),
    .Y(_01815_));
 sky130_fd_sc_hd__o2bb2ai_2 _25996_ (.A1_N(_01810_),
    .A2_N(_01811_),
    .B1(_01813_),
    .B2(_01475_),
    .Y(_01816_));
 sky130_fd_sc_hd__o2111ai_4 _25997_ (.A1(net252),
    .A2(_01471_),
    .B1(_01810_),
    .C1(_01811_),
    .D1(_01814_),
    .Y(_01817_));
 sky130_fd_sc_hd__nand3_1 _25998_ (.A(_01816_),
    .B(_01817_),
    .C(net159),
    .Y(_01818_));
 sky130_fd_sc_hd__a31o_1 _25999_ (.A1(_01816_),
    .A2(_01817_),
    .A3(net159),
    .B1(_01806_),
    .X(_01819_));
 sky130_fd_sc_hd__o311a_1 _26000_ (.A1(_05765_),
    .A2(net288),
    .A3(_01156_),
    .B1(_01165_),
    .C1(_01489_),
    .X(_01821_));
 sky130_fd_sc_hd__a22oi_1 _26001_ (.A1(_01159_),
    .A2(_01165_),
    .B1(_01487_),
    .B2(net254),
    .Y(_01822_));
 sky130_fd_sc_hd__a21o_1 _26002_ (.A1(_01490_),
    .A2(_01494_),
    .B1(_01488_),
    .X(_01823_));
 sky130_fd_sc_hd__a31oi_1 _26003_ (.A1(_01816_),
    .A2(_01817_),
    .A3(net159),
    .B1(net252),
    .Y(_01824_));
 sky130_fd_sc_hd__a311oi_2 _26004_ (.A1(_01816_),
    .A2(_01817_),
    .A3(net159),
    .B1(_01806_),
    .C1(net252),
    .Y(_01825_));
 sky130_fd_sc_hd__a311o_1 _26005_ (.A1(_01816_),
    .A2(_01817_),
    .A3(net159),
    .B1(_01806_),
    .C1(net252),
    .X(_01826_));
 sky130_fd_sc_hd__a2bb2oi_2 _26006_ (.A1_N(net284),
    .A2_N(net281),
    .B1(_01807_),
    .B2(_01818_),
    .Y(_01827_));
 sky130_fd_sc_hd__a22o_1 _26007_ (.A1(_06306_),
    .A2(_06308_),
    .B1(_01807_),
    .B2(_01818_),
    .X(_01828_));
 sky130_fd_sc_hd__o211ai_1 _26008_ (.A1(_01492_),
    .A2(_01821_),
    .B1(_01826_),
    .C1(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__o22ai_1 _26009_ (.A1(_01488_),
    .A2(_01822_),
    .B1(_01825_),
    .B2(_01827_),
    .Y(_01830_));
 sky130_fd_sc_hd__nand3_2 _26010_ (.A(_01829_),
    .B(_01830_),
    .C(net149),
    .Y(_01832_));
 sky130_fd_sc_hd__a22o_1 _26011_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_01807_),
    .B2(_01818_),
    .X(_01833_));
 sky130_fd_sc_hd__nand3_1 _26012_ (.A(_01828_),
    .B(_01823_),
    .C(_01826_),
    .Y(_01834_));
 sky130_fd_sc_hd__o22ai_1 _26013_ (.A1(_01492_),
    .A2(_01821_),
    .B1(_01825_),
    .B2(_01827_),
    .Y(_01835_));
 sky130_fd_sc_hd__o211ai_1 _26014_ (.A1(_08709_),
    .A2(_08712_),
    .B1(_01834_),
    .C1(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__o21ai_2 _26015_ (.A1(net149),
    .A2(_01819_),
    .B1(_01832_),
    .Y(_01837_));
 sky130_fd_sc_hd__o211a_1 _26016_ (.A1(_01819_),
    .A2(net149),
    .B1(_06014_),
    .C1(_01832_),
    .X(_01838_));
 sky130_fd_sc_hd__o211ai_2 _26017_ (.A1(_01819_),
    .A2(net149),
    .B1(_06014_),
    .C1(_01832_),
    .Y(_01839_));
 sky130_fd_sc_hd__and3_1 _26018_ (.A(_01836_),
    .B(net254),
    .C(_01833_),
    .X(_01840_));
 sky130_fd_sc_hd__o211ai_2 _26019_ (.A1(net285),
    .A2(_06012_),
    .B1(_01833_),
    .C1(_01836_),
    .Y(_01841_));
 sky130_fd_sc_hd__a21oi_1 _26020_ (.A1(_01507_),
    .A2(_01508_),
    .B1(_01500_),
    .Y(_01843_));
 sky130_fd_sc_hd__a31o_1 _26021_ (.A1(_01503_),
    .A2(_01507_),
    .A3(_01508_),
    .B1(_01500_),
    .X(_01844_));
 sky130_fd_sc_hd__o2bb2ai_1 _26022_ (.A1_N(_01839_),
    .A2_N(_01841_),
    .B1(_01843_),
    .B2(_01501_),
    .Y(_01845_));
 sky130_fd_sc_hd__nand3_1 _26023_ (.A(_01844_),
    .B(_01841_),
    .C(_01839_),
    .Y(_01846_));
 sky130_fd_sc_hd__o211ai_4 _26024_ (.A1(net148),
    .A2(net147),
    .B1(_01845_),
    .C1(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__or3_2 _26025_ (.A(net148),
    .B(net147),
    .C(_01837_),
    .X(_01848_));
 sky130_fd_sc_hd__o31a_2 _26026_ (.A1(net148),
    .A2(net147),
    .A3(_01837_),
    .B1(_01847_),
    .X(_01849_));
 sky130_fd_sc_hd__a21oi_4 _26027_ (.A1(_01847_),
    .A2(_01848_),
    .B1(net263),
    .Y(_01850_));
 sky130_fd_sc_hd__o221a_1 _26028_ (.A1(_05765_),
    .A2(net288),
    .B1(net146),
    .B2(_01837_),
    .C1(_01847_),
    .X(_01851_));
 sky130_fd_sc_hd__o221ai_4 _26029_ (.A1(_05765_),
    .A2(net288),
    .B1(net146),
    .B2(_01837_),
    .C1(_01847_),
    .Y(_01852_));
 sky130_fd_sc_hd__a31oi_1 _26030_ (.A1(_04238_),
    .A2(_00821_),
    .A3(_00832_),
    .B1(_00448_),
    .Y(_01854_));
 sky130_fd_sc_hd__nand4_2 _26031_ (.A(_01193_),
    .B(_01854_),
    .C(_01196_),
    .D(_00842_),
    .Y(_01855_));
 sky130_fd_sc_hd__a31oi_4 _26032_ (.A1(_01514_),
    .A2(_01515_),
    .A3(_05507_),
    .B1(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__a31o_1 _26033_ (.A1(_01514_),
    .A2(_01515_),
    .A3(_05507_),
    .B1(_01855_),
    .X(_01857_));
 sky130_fd_sc_hd__a211oi_4 _26034_ (.A1(_01525_),
    .A2(_01521_),
    .B1(_01522_),
    .C1(_01856_),
    .Y(_01858_));
 sky130_fd_sc_hd__o211ai_4 _26035_ (.A1(_01526_),
    .A2(_01520_),
    .B1(_01523_),
    .C1(_01857_),
    .Y(_01859_));
 sky130_fd_sc_hd__o211a_1 _26036_ (.A1(_05507_),
    .A2(_01517_),
    .B1(_00459_),
    .C1(_01856_),
    .X(_01860_));
 sky130_fd_sc_hd__o211ai_4 _26037_ (.A1(_05507_),
    .A2(_01517_),
    .B1(_00459_),
    .C1(_01856_),
    .Y(_01861_));
 sky130_fd_sc_hd__a31o_1 _26038_ (.A1(_01523_),
    .A2(_01528_),
    .A3(_01857_),
    .B1(_01860_),
    .X(_01862_));
 sky130_fd_sc_hd__nand2_1 _26039_ (.A(_01852_),
    .B(_01861_),
    .Y(_01863_));
 sky130_fd_sc_hd__nand4b_4 _26040_ (.A_N(_01850_),
    .B(_01852_),
    .C(_01859_),
    .D(_01861_),
    .Y(_01865_));
 sky130_fd_sc_hd__o22ai_4 _26041_ (.A1(_01850_),
    .A2(_01851_),
    .B1(_01858_),
    .B2(_01860_),
    .Y(_01866_));
 sky130_fd_sc_hd__o211ai_4 _26042_ (.A1(_09553_),
    .A2(_09556_),
    .B1(_01865_),
    .C1(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__a21oi_1 _26043_ (.A1(_01847_),
    .A2(_01848_),
    .B1(_09563_),
    .Y(_01868_));
 sky130_fd_sc_hd__or3_2 _26044_ (.A(_09553_),
    .B(net155),
    .C(_01849_),
    .X(_01869_));
 sky130_fd_sc_hd__a31oi_4 _26045_ (.A1(_09563_),
    .A2(_01865_),
    .A3(_01866_),
    .B1(_01868_),
    .Y(_01870_));
 sky130_fd_sc_hd__a21oi_1 _26046_ (.A1(_01867_),
    .A2(_01869_),
    .B1(_09579_),
    .Y(_01871_));
 sky130_fd_sc_hd__or3_2 _26047_ (.A(net142),
    .B(_09573_),
    .C(_01870_),
    .X(_01872_));
 sky130_fd_sc_hd__a31oi_1 _26048_ (.A1(_09563_),
    .A2(_01865_),
    .A3(_01866_),
    .B1(net292),
    .Y(_01873_));
 sky130_fd_sc_hd__o211a_4 _26049_ (.A1(_09563_),
    .A2(_01849_),
    .B1(_05507_),
    .C1(_01867_),
    .X(_01874_));
 sky130_fd_sc_hd__o211ai_2 _26050_ (.A1(_09563_),
    .A2(_01849_),
    .B1(_05507_),
    .C1(_01867_),
    .Y(_01876_));
 sky130_fd_sc_hd__a21oi_4 _26051_ (.A1(_01867_),
    .A2(_01869_),
    .B1(_05507_),
    .Y(_01877_));
 sky130_fd_sc_hd__a22o_1 _26052_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_01867_),
    .B2(_01869_),
    .X(_01878_));
 sky130_fd_sc_hd__a21oi_1 _26053_ (.A1(_01869_),
    .A2(_01873_),
    .B1(_01877_),
    .Y(_01879_));
 sky130_fd_sc_hd__a21oi_4 _26054_ (.A1(_01537_),
    .A2(_01533_),
    .B1(_01538_),
    .Y(_01880_));
 sky130_fd_sc_hd__o21a_2 _26055_ (.A1(_01874_),
    .A2(_01877_),
    .B1(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__o21ai_2 _26056_ (.A1(_01874_),
    .A2(_01877_),
    .B1(_01880_),
    .Y(_01882_));
 sky130_fd_sc_hd__nand3b_2 _26057_ (.A_N(_01880_),
    .B(_01878_),
    .C(_01876_),
    .Y(_01883_));
 sky130_fd_sc_hd__o31ai_4 _26058_ (.A1(_01880_),
    .A2(_01877_),
    .A3(_01874_),
    .B1(_09579_),
    .Y(_01884_));
 sky130_fd_sc_hd__nand3_1 _26059_ (.A(_09579_),
    .B(_01882_),
    .C(_01883_),
    .Y(_01885_));
 sky130_fd_sc_hd__a31oi_4 _26060_ (.A1(_09579_),
    .A2(_01882_),
    .A3(_01883_),
    .B1(_01871_),
    .Y(_01887_));
 sky130_fd_sc_hd__o21ai_4 _26061_ (.A1(_01881_),
    .A2(_01884_),
    .B1(_01872_),
    .Y(_01888_));
 sky130_fd_sc_hd__o211a_1 _26062_ (.A1(_01226_),
    .A2(_01216_),
    .B1(_01214_),
    .C1(_01550_),
    .X(_01889_));
 sky130_fd_sc_hd__a31oi_2 _26063_ (.A1(_01214_),
    .A2(_01234_),
    .A3(_01550_),
    .B1(_01552_),
    .Y(_01890_));
 sky130_fd_sc_hd__o221a_1 _26064_ (.A1(_09579_),
    .A2(_01870_),
    .B1(_01881_),
    .B2(_01884_),
    .C1(_05248_),
    .X(_01891_));
 sky130_fd_sc_hd__o221ai_4 _26065_ (.A1(_09579_),
    .A2(_01870_),
    .B1(_01881_),
    .B2(_01884_),
    .C1(_05248_),
    .Y(_01892_));
 sky130_fd_sc_hd__a22oi_4 _26066_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_01872_),
    .B2(_01885_),
    .Y(_01893_));
 sky130_fd_sc_hd__o21ai_1 _26067_ (.A1(net318),
    .A2(net315),
    .B1(_01888_),
    .Y(_01894_));
 sky130_fd_sc_hd__nand3_1 _26068_ (.A(_01894_),
    .B(_01890_),
    .C(_01892_),
    .Y(_01895_));
 sky130_fd_sc_hd__o22ai_2 _26069_ (.A1(_01552_),
    .A2(_01889_),
    .B1(_01891_),
    .B2(_01893_),
    .Y(_01896_));
 sky130_fd_sc_hd__or3_1 _26070_ (.A(_10474_),
    .B(net138),
    .C(_01887_),
    .X(_01898_));
 sky130_fd_sc_hd__o211ai_4 _26071_ (.A1(_10474_),
    .A2(_10475_),
    .B1(_01895_),
    .C1(_01896_),
    .Y(_01899_));
 sky130_fd_sc_hd__o21ai_2 _26072_ (.A1(net131),
    .A2(_01887_),
    .B1(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__o211a_1 _26073_ (.A1(net131),
    .A2(_01887_),
    .B1(_04227_),
    .C1(_01899_),
    .X(_01901_));
 sky130_fd_sc_hd__a21oi_2 _26074_ (.A1(_01898_),
    .A2(_01899_),
    .B1(_04227_),
    .Y(_01902_));
 sky130_fd_sc_hd__a211o_1 _26075_ (.A1(_01566_),
    .A2(_01578_),
    .B1(_01901_),
    .C1(_01902_),
    .X(_01903_));
 sky130_fd_sc_hd__o221ai_4 _26076_ (.A1(_02137_),
    .A2(_01564_),
    .B1(_01901_),
    .B2(_01902_),
    .C1(_01578_),
    .Y(_01904_));
 sky130_fd_sc_hd__o211ai_4 _26077_ (.A1(_10949_),
    .A2(net136),
    .B1(_01903_),
    .C1(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__a211o_2 _26078_ (.A1(_01898_),
    .A2(_01899_),
    .B1(_10949_),
    .C1(_10951_),
    .X(_01906_));
 sky130_fd_sc_hd__a21oi_2 _26079_ (.A1(_01905_),
    .A2(_01906_),
    .B1(_02137_),
    .Y(_01907_));
 sky130_fd_sc_hd__a22o_1 _26080_ (.A1(_02060_),
    .A2(_02082_),
    .B1(_01905_),
    .B2(_01906_),
    .X(_01909_));
 sky130_fd_sc_hd__a31oi_1 _26081_ (.A1(_10954_),
    .A2(_01903_),
    .A3(_01904_),
    .B1(_02148_),
    .Y(_01910_));
 sky130_fd_sc_hd__o211ai_4 _26082_ (.A1(_02093_),
    .A2(_02115_),
    .B1(_01905_),
    .C1(_01906_),
    .Y(_01911_));
 sky130_fd_sc_hd__nor3_1 _26083_ (.A(_00507_),
    .B(_00896_),
    .C(_00897_),
    .Y(_01912_));
 sky130_fd_sc_hd__nand4_1 _26084_ (.A(_01912_),
    .B(_01583_),
    .C(_01253_),
    .D(_01251_),
    .Y(_01913_));
 sky130_fd_sc_hd__o211ai_4 _26085_ (.A1(_01586_),
    .A2(_01582_),
    .B1(_01584_),
    .C1(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor4b_1 _26086_ (.A(_00508_),
    .B(_01249_),
    .C(_01252_),
    .D_N(_01912_),
    .Y(_01915_));
 sky130_fd_sc_hd__nand3_4 _26087_ (.A(_01915_),
    .B(_01584_),
    .C(_01583_),
    .Y(_01916_));
 sky130_fd_sc_hd__nand2_2 _26088_ (.A(_01914_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__a221oi_2 _26089_ (.A1(_01906_),
    .A2(_01910_),
    .B1(_01914_),
    .B2(_01916_),
    .C1(_01907_),
    .Y(_01918_));
 sky130_fd_sc_hd__a21oi_1 _26090_ (.A1(_01909_),
    .A2(_01911_),
    .B1(_01917_),
    .Y(_01920_));
 sky130_fd_sc_hd__a211o_2 _26091_ (.A1(_01905_),
    .A2(_01906_),
    .B1(_11459_),
    .C1(_11461_),
    .X(_01921_));
 sky130_fd_sc_hd__o21ai_4 _26092_ (.A1(_01918_),
    .A2(_01920_),
    .B1(_11465_),
    .Y(_01922_));
 sky130_fd_sc_hd__and3_1 _26093_ (.A(_01922_),
    .B(_00240_),
    .C(_01921_),
    .X(_01923_));
 sky130_fd_sc_hd__o211ai_1 _26094_ (.A1(_00218_),
    .A2(_00229_),
    .B1(_01921_),
    .C1(_01922_),
    .Y(_01924_));
 sky130_fd_sc_hd__a22o_1 _26095_ (.A1(_00185_),
    .A2(_00207_),
    .B1(_01921_),
    .B2(_01922_),
    .X(_01925_));
 sky130_fd_sc_hd__o32ai_2 _26096_ (.A1(net361),
    .A2(net345),
    .A3(_01589_),
    .B1(_01591_),
    .B2(_01594_),
    .Y(_01926_));
 sky130_fd_sc_hd__a221oi_2 _26097_ (.A1(_01594_),
    .A2(_01593_),
    .B1(_01925_),
    .B2(_01924_),
    .C1(_01591_),
    .Y(_01927_));
 sky130_fd_sc_hd__o211ai_4 _26098_ (.A1(_11944_),
    .A2(_01927_),
    .B1(_01922_),
    .C1(_01921_),
    .Y(_01928_));
 sky130_fd_sc_hd__a21oi_1 _26099_ (.A1(_05119_),
    .A2(_01597_),
    .B1(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__and3_1 _26100_ (.A(_05119_),
    .B(_01597_),
    .C(_01928_),
    .X(_01931_));
 sky130_fd_sc_hd__nor2_1 _26101_ (.A(_01929_),
    .B(_01931_),
    .Y(net101));
 sky130_fd_sc_hd__o22a_1 _26102_ (.A1(_04832_),
    .A2(_04942_),
    .B1(_01597_),
    .B2(_01928_),
    .X(_01932_));
 sky130_fd_sc_hd__o311a_1 _26103_ (.A1(_03399_),
    .A2(net24),
    .A3(_10962_),
    .B1(_01603_),
    .C1(_01608_),
    .X(_01933_));
 sky130_fd_sc_hd__o211ai_1 _26104_ (.A1(_01601_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_01608_),
    .Y(_01934_));
 sky130_fd_sc_hd__and3_2 _26105_ (.A(_01934_),
    .B(_04029_),
    .C(_05234_),
    .X(_01935_));
 sky130_fd_sc_hd__or4_1 _26106_ (.A(_03986_),
    .B(_03997_),
    .C(net271),
    .D(_01933_),
    .X(_01936_));
 sky130_fd_sc_hd__o21ai_1 _26107_ (.A1(_01614_),
    .A2(_01617_),
    .B1(_01613_),
    .Y(_01937_));
 sky130_fd_sc_hd__and3_1 _26108_ (.A(_01934_),
    .B(_04029_),
    .C(_10971_),
    .X(_01938_));
 sky130_fd_sc_hd__o22a_1 _26109_ (.A1(_10965_),
    .A2(_10967_),
    .B1(_04040_),
    .B2(_01933_),
    .X(_01939_));
 sky130_fd_sc_hd__nor2_1 _26110_ (.A(_01938_),
    .B(_01939_),
    .Y(_01941_));
 sky130_fd_sc_hd__a21boi_2 _26111_ (.A1(_01613_),
    .A2(_01619_),
    .B1_N(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__nand2_1 _26112_ (.A(_01937_),
    .B(_01941_),
    .Y(_01943_));
 sky130_fd_sc_hd__o211ai_4 _26113_ (.A1(_01938_),
    .A2(_01939_),
    .B1(_01613_),
    .C1(_01619_),
    .Y(_01944_));
 sky130_fd_sc_hd__nand3_1 _26114_ (.A(_01943_),
    .B(_01944_),
    .C(net271),
    .Y(_01945_));
 sky130_fd_sc_hd__a31oi_4 _26115_ (.A1(_01943_),
    .A2(_01944_),
    .A3(net271),
    .B1(_01935_),
    .Y(_01946_));
 sky130_fd_sc_hd__a2bb2oi_1 _26116_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_01936_),
    .B2(_01945_),
    .Y(_01947_));
 sky130_fd_sc_hd__a2bb2o_1 _26117_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_01936_),
    .B2(_01945_),
    .X(_01948_));
 sky130_fd_sc_hd__a31o_2 _26118_ (.A1(_01943_),
    .A2(_01944_),
    .A3(net271),
    .B1(_10492_),
    .X(_01949_));
 sky130_fd_sc_hd__o311a_1 _26119_ (.A1(_04040_),
    .A2(net271),
    .A3(_01933_),
    .B1(net150),
    .C1(_01945_),
    .X(_01950_));
 sky130_fd_sc_hd__nand3_1 _26120_ (.A(_01630_),
    .B(_01634_),
    .C(_01638_),
    .Y(_01952_));
 sky130_fd_sc_hd__o2bb2ai_1 _26121_ (.A1_N(_01630_),
    .A2_N(_01634_),
    .B1(net153),
    .B2(_01625_),
    .Y(_01953_));
 sky130_fd_sc_hd__a31oi_4 _26122_ (.A1(_01630_),
    .A2(_01634_),
    .A3(_01638_),
    .B1(_01639_),
    .Y(_01954_));
 sky130_fd_sc_hd__o21ai_2 _26123_ (.A1(_01947_),
    .A2(_01950_),
    .B1(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__o2111ai_4 _26124_ (.A1(_01949_),
    .A2(_01935_),
    .B1(_01638_),
    .C1(_01948_),
    .D1(_01953_),
    .Y(_01956_));
 sky130_fd_sc_hd__a2bb2o_2 _26125_ (.A1_N(_05478_),
    .A2_N(_05479_),
    .B1(_01936_),
    .B2(_01945_),
    .X(_01957_));
 sky130_fd_sc_hd__inv_2 _26126_ (.A(_01957_),
    .Y(_01958_));
 sky130_fd_sc_hd__o311a_1 _26127_ (.A1(_01947_),
    .A2(_01950_),
    .A3(_01954_),
    .B1(net244),
    .C1(_01955_),
    .X(_01959_));
 sky130_fd_sc_hd__nand3_2 _26128_ (.A(_01956_),
    .B(net244),
    .C(_01955_),
    .Y(_01960_));
 sky130_fd_sc_hd__a31o_2 _26129_ (.A1(_01956_),
    .A2(net244),
    .A3(_01955_),
    .B1(_01958_),
    .X(_01961_));
 sky130_fd_sc_hd__o31a_1 _26130_ (.A1(net270),
    .A2(net268),
    .A3(_01946_),
    .B1(_01960_),
    .X(_01963_));
 sky130_fd_sc_hd__a2bb2oi_2 _26131_ (.A1_N(net170),
    .A2_N(_10022_),
    .B1(_01957_),
    .B2(_01960_),
    .Y(_01964_));
 sky130_fd_sc_hd__o22ai_4 _26132_ (.A1(net170),
    .A2(net168),
    .B1(_01958_),
    .B2(_01959_),
    .Y(_01965_));
 sky130_fd_sc_hd__a31oi_1 _26133_ (.A1(_01956_),
    .A2(net244),
    .A3(_01955_),
    .B1(net151),
    .Y(_01966_));
 sky130_fd_sc_hd__o211ai_4 _26134_ (.A1(net244),
    .A2(_01946_),
    .B1(net153),
    .C1(_01960_),
    .Y(_01967_));
 sky130_fd_sc_hd__a21oi_1 _26135_ (.A1(_01957_),
    .A2(_01966_),
    .B1(_01964_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _26136_ (.A(_01965_),
    .B(_01967_),
    .Y(_01969_));
 sky130_fd_sc_hd__and3_1 _26137_ (.A(_00623_),
    .B(_00994_),
    .C(_00995_),
    .X(_01970_));
 sky130_fd_sc_hd__nor4_1 _26138_ (.A(_00625_),
    .B(_00996_),
    .C(_01340_),
    .D(_01342_),
    .Y(_01971_));
 sky130_fd_sc_hd__nand3_1 _26139_ (.A(_01656_),
    .B(_01970_),
    .C(_01344_),
    .Y(_01972_));
 sky130_fd_sc_hd__o211ai_4 _26140_ (.A1(_01660_),
    .A2(_01654_),
    .B1(_01657_),
    .C1(_01972_),
    .Y(_01974_));
 sky130_fd_sc_hd__nand4b_4 _26141_ (.A_N(_00636_),
    .B(_01656_),
    .C(_01971_),
    .D(_01657_),
    .Y(_01975_));
 sky130_fd_sc_hd__nand2_1 _26142_ (.A(_01974_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__a21oi_1 _26143_ (.A1(_01974_),
    .A2(_01975_),
    .B1(_01969_),
    .Y(_01977_));
 sky130_fd_sc_hd__o22ai_2 _26144_ (.A1(net265),
    .A2(net264),
    .B1(_01968_),
    .B2(_01976_),
    .Y(_01978_));
 sky130_fd_sc_hd__nand4_4 _26145_ (.A(_01965_),
    .B(_01967_),
    .C(_01974_),
    .D(_01975_),
    .Y(_01979_));
 sky130_fd_sc_hd__a22o_1 _26146_ (.A1(_01965_),
    .A2(_01967_),
    .B1(_01974_),
    .B2(_01975_),
    .X(_01980_));
 sky130_fd_sc_hd__a21oi_2 _26147_ (.A1(_01957_),
    .A2(_01960_),
    .B1(_05752_),
    .Y(_01981_));
 sky130_fd_sc_hd__or3_2 _26148_ (.A(net265),
    .B(net264),
    .C(_01963_),
    .X(_01982_));
 sky130_fd_sc_hd__nand3_2 _26149_ (.A(_01980_),
    .B(_05752_),
    .C(_01979_),
    .Y(_01983_));
 sky130_fd_sc_hd__a31o_2 _26150_ (.A1(_01980_),
    .A2(_05752_),
    .A3(_01979_),
    .B1(_01981_),
    .X(_01985_));
 sky130_fd_sc_hd__a211o_1 _26151_ (.A1(_01982_),
    .A2(_01983_),
    .B1(net260),
    .C1(net255),
    .X(_01986_));
 sky130_fd_sc_hd__a311oi_4 _26152_ (.A1(_01980_),
    .A2(_05752_),
    .A3(_01979_),
    .B1(_01981_),
    .C1(net171),
    .Y(_01987_));
 sky130_fd_sc_hd__nand3_4 _26153_ (.A(_01983_),
    .B(net172),
    .C(_01982_),
    .Y(_01988_));
 sky130_fd_sc_hd__o221ai_4 _26154_ (.A1(_05752_),
    .A2(_01961_),
    .B1(_01977_),
    .B2(_01978_),
    .C1(net171),
    .Y(_01989_));
 sky130_fd_sc_hd__o221a_1 _26155_ (.A1(_01353_),
    .A2(net177),
    .B1(net174),
    .B2(_01668_),
    .C1(_01671_),
    .X(_01990_));
 sky130_fd_sc_hd__o211ai_1 _26156_ (.A1(_08731_),
    .A2(_01352_),
    .B1(_01670_),
    .C1(_01674_),
    .Y(_01991_));
 sky130_fd_sc_hd__o21ai_2 _26157_ (.A1(net174),
    .A2(_01668_),
    .B1(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__a31oi_4 _26158_ (.A1(_01355_),
    .A2(_01670_),
    .A3(_01674_),
    .B1(_01675_),
    .Y(_01993_));
 sky130_fd_sc_hd__o2bb2ai_4 _26159_ (.A1_N(_01988_),
    .A2_N(_01989_),
    .B1(_01990_),
    .B2(_01673_),
    .Y(_01994_));
 sky130_fd_sc_hd__nand3_1 _26160_ (.A(_01988_),
    .B(_01989_),
    .C(_01992_),
    .Y(_01996_));
 sky130_fd_sc_hd__a31oi_4 _26161_ (.A1(_01988_),
    .A2(_01989_),
    .A3(_01992_),
    .B1(_05995_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand3_1 _26162_ (.A(net240),
    .B(_01994_),
    .C(_01996_),
    .Y(_01998_));
 sky130_fd_sc_hd__a22oi_4 _26163_ (.A1(_05995_),
    .A2(_01985_),
    .B1(_01997_),
    .B2(_01994_),
    .Y(_01999_));
 sky130_fd_sc_hd__a22o_1 _26164_ (.A1(_05995_),
    .A2(_01985_),
    .B1(_01997_),
    .B2(_01994_),
    .X(_02000_));
 sky130_fd_sc_hd__o221a_1 _26165_ (.A1(net200),
    .A2(_01368_),
    .B1(_01694_),
    .B2(_01383_),
    .C1(_01690_),
    .X(_02001_));
 sky130_fd_sc_hd__o221ai_2 _26166_ (.A1(net200),
    .A2(_01368_),
    .B1(_01694_),
    .B2(_01383_),
    .C1(_01690_),
    .Y(_02002_));
 sky130_fd_sc_hd__a2bb2oi_1 _26167_ (.A1_N(_01686_),
    .A2_N(_08731_),
    .B1(_01373_),
    .B2(_01695_),
    .Y(_02003_));
 sky130_fd_sc_hd__a21oi_1 _26168_ (.A1(_01997_),
    .A2(_01994_),
    .B1(net173),
    .Y(_02004_));
 sky130_fd_sc_hd__a221oi_2 _26169_ (.A1(_05995_),
    .A2(_01985_),
    .B1(_01997_),
    .B2(_01994_),
    .C1(net173),
    .Y(_02005_));
 sky130_fd_sc_hd__nand3_1 _26170_ (.A(_01998_),
    .B(net174),
    .C(_01986_),
    .Y(_02007_));
 sky130_fd_sc_hd__a2bb2oi_2 _26171_ (.A1_N(net194),
    .A2_N(net192),
    .B1(_01986_),
    .B2(_01998_),
    .Y(_02008_));
 sky130_fd_sc_hd__a2bb2o_1 _26172_ (.A1_N(net194),
    .A2_N(net192),
    .B1(_01986_),
    .B2(_01998_),
    .X(_02009_));
 sky130_fd_sc_hd__o211ai_1 _26173_ (.A1(_01691_),
    .A2(_02001_),
    .B1(_02007_),
    .C1(_02009_),
    .Y(_02010_));
 sky130_fd_sc_hd__o22ai_1 _26174_ (.A1(_01689_),
    .A2(_02003_),
    .B1(_02005_),
    .B2(_02008_),
    .Y(_02011_));
 sky130_fd_sc_hd__nand3_1 _26175_ (.A(_02010_),
    .B(_02011_),
    .C(_06293_),
    .Y(_02012_));
 sky130_fd_sc_hd__o211ai_1 _26176_ (.A1(_01689_),
    .A2(_02003_),
    .B1(_02007_),
    .C1(_02009_),
    .Y(_02013_));
 sky130_fd_sc_hd__o22ai_1 _26177_ (.A1(_01691_),
    .A2(_02001_),
    .B1(_02005_),
    .B2(_02008_),
    .Y(_02014_));
 sky130_fd_sc_hd__nand3_2 _26178_ (.A(_02013_),
    .B(_02014_),
    .C(_06293_),
    .Y(_02015_));
 sky130_fd_sc_hd__o31a_2 _26179_ (.A1(net239),
    .A2(_06292_),
    .A3(_01999_),
    .B1(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__o211ai_4 _26180_ (.A1(_02000_),
    .A2(_06293_),
    .B1(_08731_),
    .C1(_02012_),
    .Y(_02017_));
 sky130_fd_sc_hd__o211a_1 _26181_ (.A1(_06293_),
    .A2(_01999_),
    .B1(net178),
    .C1(_02015_),
    .X(_02018_));
 sky130_fd_sc_hd__o211ai_4 _26182_ (.A1(_06293_),
    .A2(_01999_),
    .B1(net178),
    .C1(_02015_),
    .Y(_02019_));
 sky130_fd_sc_hd__nand2_1 _26183_ (.A(_02017_),
    .B(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__o2bb2ai_2 _26184_ (.A1_N(_01724_),
    .A2_N(_01726_),
    .B1(net200),
    .B2(_01707_),
    .Y(_02021_));
 sky130_fd_sc_hd__nand2_1 _26185_ (.A(_01713_),
    .B(_01726_),
    .Y(_02022_));
 sky130_fd_sc_hd__a31oi_4 _26186_ (.A1(_01713_),
    .A2(_01724_),
    .A3(_01726_),
    .B1(_01709_),
    .Y(_02023_));
 sky130_fd_sc_hd__o2111ai_1 _26187_ (.A1(_08314_),
    .A2(_01708_),
    .B1(_02017_),
    .C1(_02019_),
    .D1(_02021_),
    .Y(_02024_));
 sky130_fd_sc_hd__a22oi_4 _26188_ (.A1(_02017_),
    .A2(_02019_),
    .B1(_02021_),
    .B2(_01713_),
    .Y(_02025_));
 sky130_fd_sc_hd__o221ai_1 _26189_ (.A1(net200),
    .A2(_01707_),
    .B1(_01715_),
    .B2(_01728_),
    .C1(_02020_),
    .Y(_02026_));
 sky130_fd_sc_hd__o22ai_4 _26190_ (.A1(net238),
    .A2(net236),
    .B1(_02020_),
    .B2(_02023_),
    .Y(_02028_));
 sky130_fd_sc_hd__nand3_1 _26191_ (.A(_02024_),
    .B(_02026_),
    .C(net209),
    .Y(_02029_));
 sky130_fd_sc_hd__or3_1 _26192_ (.A(net238),
    .B(net236),
    .C(_02016_),
    .X(_02030_));
 sky130_fd_sc_hd__o32a_1 _26193_ (.A1(net238),
    .A2(net236),
    .A3(_02016_),
    .B1(_02025_),
    .B2(_02028_),
    .X(_02031_));
 sky130_fd_sc_hd__o22ai_4 _26194_ (.A1(net209),
    .A2(_02016_),
    .B1(_02025_),
    .B2(_02028_),
    .Y(_02032_));
 sky130_fd_sc_hd__a22oi_4 _26195_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_02029_),
    .B2(_02030_),
    .Y(_02033_));
 sky130_fd_sc_hd__o21ai_4 _26196_ (.A1(_08307_),
    .A2(net216),
    .B1(_02032_),
    .Y(_02034_));
 sky130_fd_sc_hd__o22a_1 _26197_ (.A1(_08311_),
    .A2(net215),
    .B1(_02025_),
    .B2(_02028_),
    .X(_02035_));
 sky130_fd_sc_hd__o221ai_4 _26198_ (.A1(net209),
    .A2(_02016_),
    .B1(_02025_),
    .B2(_02028_),
    .C1(net200),
    .Y(_02036_));
 sky130_fd_sc_hd__a21oi_1 _26199_ (.A1(_02030_),
    .A2(_02035_),
    .B1(_02033_),
    .Y(_02037_));
 sky130_fd_sc_hd__nand2_1 _26200_ (.A(_02034_),
    .B(_02036_),
    .Y(_02039_));
 sky130_fd_sc_hd__and3_1 _26201_ (.A(_00702_),
    .B(_01068_),
    .C(_01070_),
    .X(_02040_));
 sky130_fd_sc_hd__nor3b_1 _26202_ (.A(_01412_),
    .B(_01415_),
    .C_N(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand3_1 _26203_ (.A(_01740_),
    .B(_02040_),
    .C(_01417_),
    .Y(_02042_));
 sky130_fd_sc_hd__o211ai_4 _26204_ (.A1(_01745_),
    .A2(_01739_),
    .B1(_01741_),
    .C1(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__inv_2 _26205_ (.A(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__nand3_1 _26206_ (.A(_02041_),
    .B(_01741_),
    .C(_00710_),
    .Y(_02045_));
 sky130_fd_sc_hd__nand4_4 _26207_ (.A(_02041_),
    .B(_01741_),
    .C(_01740_),
    .D(_00710_),
    .Y(_02046_));
 sky130_fd_sc_hd__inv_2 _26208_ (.A(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__o21ai_1 _26209_ (.A1(_01739_),
    .A2(_02045_),
    .B1(_02043_),
    .Y(_02048_));
 sky130_fd_sc_hd__a21oi_2 _26210_ (.A1(_02043_),
    .A2(_02046_),
    .B1(_02039_),
    .Y(_02050_));
 sky130_fd_sc_hd__o22ai_2 _26211_ (.A1(net229),
    .A2(net228),
    .B1(_02037_),
    .B2(_02048_),
    .Y(_02051_));
 sky130_fd_sc_hd__and3_1 _26212_ (.A(_06900_),
    .B(_06902_),
    .C(_02032_),
    .X(_02052_));
 sky130_fd_sc_hd__or3_1 _26213_ (.A(net229),
    .B(net228),
    .C(_02031_),
    .X(_02053_));
 sky130_fd_sc_hd__nand4_2 _26214_ (.A(_02034_),
    .B(_02036_),
    .C(_02043_),
    .D(_02046_),
    .Y(_02054_));
 sky130_fd_sc_hd__a22o_1 _26215_ (.A1(_02034_),
    .A2(_02036_),
    .B1(_02043_),
    .B2(_02046_),
    .X(_02055_));
 sky130_fd_sc_hd__nand3_2 _26216_ (.A(_02055_),
    .B(_06903_),
    .C(_02054_),
    .Y(_02056_));
 sky130_fd_sc_hd__a31o_1 _26217_ (.A1(_02055_),
    .A2(_06903_),
    .A3(_02054_),
    .B1(_02052_),
    .X(_02057_));
 sky130_fd_sc_hd__o221a_1 _26218_ (.A1(_06903_),
    .A2(_02032_),
    .B1(_02050_),
    .B2(_02051_),
    .C1(_07232_),
    .X(_02058_));
 sky130_fd_sc_hd__a211o_2 _26219_ (.A1(_02053_),
    .A2(_02056_),
    .B1(net207),
    .C1(net205),
    .X(_02059_));
 sky130_fd_sc_hd__a311oi_2 _26220_ (.A1(_02055_),
    .A2(_06903_),
    .A3(_02054_),
    .B1(_07936_),
    .C1(_02052_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand3_4 _26221_ (.A(_02056_),
    .B(_07935_),
    .C(_02053_),
    .Y(_02062_));
 sky130_fd_sc_hd__o221ai_4 _26222_ (.A1(_06903_),
    .A2(_02032_),
    .B1(_02050_),
    .B2(_02051_),
    .C1(_07936_),
    .Y(_02063_));
 sky130_fd_sc_hd__a21oi_1 _26223_ (.A1(_01428_),
    .A2(_01758_),
    .B1(_01755_),
    .Y(_02064_));
 sky130_fd_sc_hd__o221a_1 _26224_ (.A1(_01423_),
    .A2(net223),
    .B1(net202),
    .B2(_01749_),
    .C1(_01758_),
    .X(_02065_));
 sky130_fd_sc_hd__a31oi_2 _26225_ (.A1(_01428_),
    .A2(_01753_),
    .A3(_01758_),
    .B1(_01755_),
    .Y(_02066_));
 sky130_fd_sc_hd__a21boi_1 _26226_ (.A1(_02062_),
    .A2(_02063_),
    .B1_N(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__o2bb2ai_2 _26227_ (.A1_N(_02062_),
    .A2_N(_02063_),
    .B1(_02064_),
    .B2(_01752_),
    .Y(_02068_));
 sky130_fd_sc_hd__o211a_1 _26228_ (.A1(_01755_),
    .A2(_02065_),
    .B1(_02063_),
    .C1(_02062_),
    .X(_02069_));
 sky130_fd_sc_hd__o211ai_4 _26229_ (.A1(_01755_),
    .A2(_02065_),
    .B1(_02063_),
    .C1(_02062_),
    .Y(_02070_));
 sky130_fd_sc_hd__o211ai_4 _26230_ (.A1(net207),
    .A2(net205),
    .B1(_02068_),
    .C1(_02070_),
    .Y(_02072_));
 sky130_fd_sc_hd__o22ai_2 _26231_ (.A1(net207),
    .A2(net205),
    .B1(_02067_),
    .B2(_02069_),
    .Y(_02073_));
 sky130_fd_sc_hd__o31a_1 _26232_ (.A1(_07232_),
    .A2(_02067_),
    .A3(_02069_),
    .B1(_02059_),
    .X(_02074_));
 sky130_fd_sc_hd__a31o_2 _26233_ (.A1(_07233_),
    .A2(_02068_),
    .A3(_02070_),
    .B1(_02058_),
    .X(_02075_));
 sky130_fd_sc_hd__o221ai_4 _26234_ (.A1(_06922_),
    .A2(_01435_),
    .B1(_07246_),
    .B2(_01767_),
    .C1(_01449_),
    .Y(_02076_));
 sky130_fd_sc_hd__a31oi_1 _26235_ (.A1(_01437_),
    .A2(_01449_),
    .A3(_01768_),
    .B1(_01769_),
    .Y(_02077_));
 sky130_fd_sc_hd__a31o_1 _26236_ (.A1(_07233_),
    .A2(_02068_),
    .A3(_02070_),
    .B1(net202),
    .X(_02078_));
 sky130_fd_sc_hd__a311oi_1 _26237_ (.A1(_07233_),
    .A2(_02068_),
    .A3(_02070_),
    .B1(net202),
    .C1(_02058_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand3_4 _26238_ (.A(_02072_),
    .B(_07564_),
    .C(_02059_),
    .Y(_02080_));
 sky130_fd_sc_hd__a22oi_4 _26239_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_02059_),
    .B2(_02072_),
    .Y(_02081_));
 sky130_fd_sc_hd__o221ai_4 _26240_ (.A1(net221),
    .A2(net220),
    .B1(_02057_),
    .B2(_07233_),
    .C1(_02073_),
    .Y(_02083_));
 sky130_fd_sc_hd__o2111ai_4 _26241_ (.A1(_01769_),
    .A2(_01773_),
    .B1(_02080_),
    .C1(_02083_),
    .D1(_01768_),
    .Y(_02084_));
 sky130_fd_sc_hd__o21ai_1 _26242_ (.A1(_02079_),
    .A2(_02081_),
    .B1(_02077_),
    .Y(_02085_));
 sky130_fd_sc_hd__o211ai_4 _26243_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_02084_),
    .C1(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__o211ai_1 _26244_ (.A1(_02058_),
    .A2(_02078_),
    .B1(_02083_),
    .C1(_02077_),
    .Y(_02087_));
 sky130_fd_sc_hd__o2bb2ai_1 _26245_ (.A1_N(_01770_),
    .A2_N(_02076_),
    .B1(_02079_),
    .B2(_02081_),
    .Y(_02088_));
 sky130_fd_sc_hd__nand3_1 _26246_ (.A(_02087_),
    .B(_02088_),
    .C(_07548_),
    .Y(_02089_));
 sky130_fd_sc_hd__o21ai_1 _26247_ (.A1(_07548_),
    .A2(_02074_),
    .B1(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__o21ai_4 _26248_ (.A1(_07548_),
    .A2(_02075_),
    .B1(_02086_),
    .Y(_02091_));
 sky130_fd_sc_hd__o211ai_4 _26249_ (.A1(_02075_),
    .A2(_07548_),
    .B1(net223),
    .C1(_02086_),
    .Y(_02092_));
 sky130_fd_sc_hd__o211a_2 _26250_ (.A1(_07548_),
    .A2(_02074_),
    .B1(_07246_),
    .C1(_02089_),
    .X(_02094_));
 sky130_fd_sc_hd__o211ai_2 _26251_ (.A1(_07548_),
    .A2(_02074_),
    .B1(_07246_),
    .C1(_02089_),
    .Y(_02095_));
 sky130_fd_sc_hd__nand2_1 _26252_ (.A(_02092_),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__a31oi_2 _26253_ (.A1(_01786_),
    .A2(_01793_),
    .A3(_01794_),
    .B1(_01783_),
    .Y(_02097_));
 sky130_fd_sc_hd__o311a_2 _26254_ (.A1(_06918_),
    .A2(net249),
    .A3(_01781_),
    .B1(_01803_),
    .C1(_02096_),
    .X(_02098_));
 sky130_fd_sc_hd__o22ai_4 _26255_ (.A1(net183),
    .A2(net182),
    .B1(_02096_),
    .B2(_02097_),
    .Y(_02099_));
 sky130_fd_sc_hd__o22ai_4 _26256_ (.A1(net162),
    .A2(_02091_),
    .B1(_02098_),
    .B2(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__inv_2 _26257_ (.A(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__and3_4 _26258_ (.A(_08297_),
    .B(_08299_),
    .C(_02100_),
    .X(_02102_));
 sky130_fd_sc_hd__or3_1 _26259_ (.A(net181),
    .B(net179),
    .C(_02101_),
    .X(_02103_));
 sky130_fd_sc_hd__o21a_1 _26260_ (.A1(_06914_),
    .A2(net250),
    .B1(_02100_),
    .X(_02105_));
 sky130_fd_sc_hd__o21ai_4 _26261_ (.A1(_06914_),
    .A2(net250),
    .B1(_02100_),
    .Y(_02106_));
 sky130_fd_sc_hd__o221ai_4 _26262_ (.A1(net162),
    .A2(_02091_),
    .B1(_02098_),
    .B2(_02099_),
    .C1(_06922_),
    .Y(_02107_));
 sky130_fd_sc_hd__and3_1 _26263_ (.A(_01141_),
    .B(_01143_),
    .C(_00780_),
    .X(_02108_));
 sky130_fd_sc_hd__a21boi_1 _26264_ (.A1(net252),
    .A2(_01471_),
    .B1_N(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__o211ai_2 _26265_ (.A1(net252),
    .A2(_01471_),
    .B1(_02109_),
    .C1(_01810_),
    .Y(_02110_));
 sky130_fd_sc_hd__o211a_1 _26266_ (.A1(_01815_),
    .A2(_01808_),
    .B1(_01811_),
    .C1(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__o211ai_4 _26267_ (.A1(_01815_),
    .A2(_01808_),
    .B1(_01811_),
    .C1(_02110_),
    .Y(_02112_));
 sky130_fd_sc_hd__nand4_2 _26268_ (.A(_01478_),
    .B(_01144_),
    .C(_00792_),
    .D(_01476_),
    .Y(_02113_));
 sky130_fd_sc_hd__nand3b_4 _26269_ (.A_N(_02113_),
    .B(_01811_),
    .C(_01810_),
    .Y(_02114_));
 sky130_fd_sc_hd__o21ai_1 _26270_ (.A1(_01812_),
    .A2(_02113_),
    .B1(_02112_),
    .Y(_02116_));
 sky130_fd_sc_hd__a22oi_2 _26271_ (.A1(_02106_),
    .A2(_02107_),
    .B1(_02112_),
    .B2(_02114_),
    .Y(_02117_));
 sky130_fd_sc_hd__a22o_2 _26272_ (.A1(_02106_),
    .A2(_02107_),
    .B1(_02112_),
    .B2(_02114_),
    .X(_02118_));
 sky130_fd_sc_hd__o22a_2 _26273_ (.A1(net226),
    .A2(_02100_),
    .B1(_02113_),
    .B2(_01812_),
    .X(_02119_));
 sky130_fd_sc_hd__o21ai_1 _26274_ (.A1(net226),
    .A2(_02100_),
    .B1(_02114_),
    .Y(_02120_));
 sky130_fd_sc_hd__nand3_2 _26275_ (.A(_02107_),
    .B(_02112_),
    .C(_02114_),
    .Y(_02121_));
 sky130_fd_sc_hd__o2111ai_4 _26276_ (.A1(net226),
    .A2(_02100_),
    .B1(_02106_),
    .C1(_02112_),
    .D1(_02114_),
    .Y(_02122_));
 sky130_fd_sc_hd__a311oi_4 _26277_ (.A1(_02106_),
    .A2(_02119_),
    .A3(_02112_),
    .B1(_08301_),
    .C1(_02117_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand3_1 _26278_ (.A(_02118_),
    .B(_02122_),
    .C(net159),
    .Y(_02124_));
 sky130_fd_sc_hd__a31oi_4 _26279_ (.A1(_02118_),
    .A2(_02122_),
    .A3(net159),
    .B1(_02102_),
    .Y(_02125_));
 sky130_fd_sc_hd__o22a_1 _26280_ (.A1(_08705_),
    .A2(_08707_),
    .B1(_02102_),
    .B2(_02123_),
    .X(_02127_));
 sky130_fd_sc_hd__or3_2 _26281_ (.A(net157),
    .B(_08712_),
    .C(_02125_),
    .X(_02128_));
 sky130_fd_sc_hd__a31o_1 _26282_ (.A1(_02118_),
    .A2(_02122_),
    .A3(net159),
    .B1(net233),
    .X(_02129_));
 sky130_fd_sc_hd__a311oi_4 _26283_ (.A1(_02118_),
    .A2(_02122_),
    .A3(net159),
    .B1(_02102_),
    .C1(net233),
    .Y(_02130_));
 sky130_fd_sc_hd__nand3_2 _26284_ (.A(_02124_),
    .B(net235),
    .C(_02103_),
    .Y(_02131_));
 sky130_fd_sc_hd__a2bb2oi_1 _26285_ (.A1_N(_06622_),
    .A2_N(_06624_),
    .B1(_02103_),
    .B2(_02124_),
    .Y(_02132_));
 sky130_fd_sc_hd__o22ai_4 _26286_ (.A1(_06622_),
    .A2(_06624_),
    .B1(_02102_),
    .B2(_02123_),
    .Y(_02133_));
 sky130_fd_sc_hd__o32a_1 _26287_ (.A1(net284),
    .A2(net281),
    .A3(_01819_),
    .B1(_01823_),
    .B2(_01827_),
    .X(_02134_));
 sky130_fd_sc_hd__a21oi_2 _26288_ (.A1(_01826_),
    .A2(_01823_),
    .B1(_01827_),
    .Y(_02135_));
 sky130_fd_sc_hd__o21a_2 _26289_ (.A1(_02130_),
    .A2(_02132_),
    .B1(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__o21ai_2 _26290_ (.A1(_02130_),
    .A2(_02132_),
    .B1(_02135_),
    .Y(_02138_));
 sky130_fd_sc_hd__o21ai_2 _26291_ (.A1(net235),
    .A2(_02125_),
    .B1(_02134_),
    .Y(_02139_));
 sky130_fd_sc_hd__o211ai_2 _26292_ (.A1(_02102_),
    .A2(_02129_),
    .B1(_02134_),
    .C1(_02133_),
    .Y(_02140_));
 sky130_fd_sc_hd__o22ai_4 _26293_ (.A1(net157),
    .A2(_08712_),
    .B1(_02130_),
    .B2(_02139_),
    .Y(_02141_));
 sky130_fd_sc_hd__o211ai_4 _26294_ (.A1(_02130_),
    .A2(_02139_),
    .B1(net149),
    .C1(_02138_),
    .Y(_02142_));
 sky130_fd_sc_hd__o22ai_4 _26295_ (.A1(net149),
    .A2(_02125_),
    .B1(_02136_),
    .B2(_02141_),
    .Y(_02143_));
 sky130_fd_sc_hd__o311a_1 _26296_ (.A1(_05765_),
    .A2(net288),
    .A3(_01499_),
    .B1(_01511_),
    .C1(_01839_),
    .X(_02144_));
 sky130_fd_sc_hd__a21o_1 _26297_ (.A1(_01844_),
    .A2(_01841_),
    .B1(_01838_),
    .X(_02145_));
 sky130_fd_sc_hd__a21oi_1 _26298_ (.A1(_01844_),
    .A2(_01841_),
    .B1(_01838_),
    .Y(_02146_));
 sky130_fd_sc_hd__a311oi_4 _26299_ (.A1(_02138_),
    .A2(_02140_),
    .A3(net149),
    .B1(_02127_),
    .C1(net252),
    .Y(_02147_));
 sky130_fd_sc_hd__o221ai_4 _26300_ (.A1(net149),
    .A2(_02125_),
    .B1(_02136_),
    .B2(_02141_),
    .C1(_06314_),
    .Y(_02149_));
 sky130_fd_sc_hd__a2bb2oi_2 _26301_ (.A1_N(net284),
    .A2_N(net281),
    .B1(_02128_),
    .B2(_02142_),
    .Y(_02150_));
 sky130_fd_sc_hd__o21ai_2 _26302_ (.A1(net284),
    .A2(net281),
    .B1(_02143_),
    .Y(_02151_));
 sky130_fd_sc_hd__o211ai_1 _26303_ (.A1(_01840_),
    .A2(_02144_),
    .B1(_02149_),
    .C1(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__o21ai_1 _26304_ (.A1(_02147_),
    .A2(_02150_),
    .B1(_02145_),
    .Y(_02153_));
 sky130_fd_sc_hd__o211ai_2 _26305_ (.A1(net148),
    .A2(net147),
    .B1(_02152_),
    .C1(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__a21oi_2 _26306_ (.A1(_02128_),
    .A2(_02142_),
    .B1(net146),
    .Y(_02155_));
 sky130_fd_sc_hd__a211o_2 _26307_ (.A1(_02128_),
    .A2(_02142_),
    .B1(net148),
    .C1(net147),
    .X(_02156_));
 sky130_fd_sc_hd__nand3_2 _26308_ (.A(_02151_),
    .B(_02145_),
    .C(_02149_),
    .Y(_02157_));
 sky130_fd_sc_hd__o22ai_4 _26309_ (.A1(_01840_),
    .A2(_02144_),
    .B1(_02147_),
    .B2(_02150_),
    .Y(_02158_));
 sky130_fd_sc_hd__o211ai_4 _26310_ (.A1(net148),
    .A2(net147),
    .B1(_02157_),
    .C1(_02158_),
    .Y(_02160_));
 sky130_fd_sc_hd__a31o_1 _26311_ (.A1(net146),
    .A2(_02157_),
    .A3(_02158_),
    .B1(_02155_),
    .X(_02161_));
 sky130_fd_sc_hd__o211ai_4 _26312_ (.A1(net146),
    .A2(_02143_),
    .B1(_02154_),
    .C1(_06014_),
    .Y(_02162_));
 sky130_fd_sc_hd__o21ai_2 _26313_ (.A1(net285),
    .A2(_06012_),
    .B1(_02160_),
    .Y(_02163_));
 sky130_fd_sc_hd__and3_1 _26314_ (.A(_02160_),
    .B(_06013_),
    .C(_02156_),
    .X(_02164_));
 sky130_fd_sc_hd__o211ai_4 _26315_ (.A1(net285),
    .A2(_06012_),
    .B1(_02156_),
    .C1(_02160_),
    .Y(_02165_));
 sky130_fd_sc_hd__o22a_1 _26316_ (.A1(net263),
    .A2(_01849_),
    .B1(_01858_),
    .B2(_01860_),
    .X(_02166_));
 sky130_fd_sc_hd__a31oi_4 _26317_ (.A1(_01852_),
    .A2(_01859_),
    .A3(_01861_),
    .B1(_01850_),
    .Y(_02167_));
 sky130_fd_sc_hd__o22ai_4 _26318_ (.A1(net263),
    .A2(_01849_),
    .B1(_01858_),
    .B2(_01863_),
    .Y(_02168_));
 sky130_fd_sc_hd__a21oi_4 _26319_ (.A1(_02162_),
    .A2(_02165_),
    .B1(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__o2bb2ai_1 _26320_ (.A1_N(_02162_),
    .A2_N(_02165_),
    .B1(_02166_),
    .B2(_01851_),
    .Y(_02171_));
 sky130_fd_sc_hd__o211a_1 _26321_ (.A1(_02155_),
    .A2(_02163_),
    .B1(_02168_),
    .C1(_02162_),
    .X(_02172_));
 sky130_fd_sc_hd__o211ai_2 _26322_ (.A1(_02155_),
    .A2(_02163_),
    .B1(_02168_),
    .C1(_02162_),
    .Y(_02173_));
 sky130_fd_sc_hd__o22ai_2 _26323_ (.A1(net156),
    .A2(_09556_),
    .B1(_02169_),
    .B2(_02172_),
    .Y(_02174_));
 sky130_fd_sc_hd__and3_1 _26324_ (.A(_02161_),
    .B(_09557_),
    .C(_09554_),
    .X(_02175_));
 sky130_fd_sc_hd__a211o_2 _26325_ (.A1(_02156_),
    .A2(_02160_),
    .B1(net156),
    .C1(_09556_),
    .X(_02176_));
 sky130_fd_sc_hd__a31o_1 _26326_ (.A1(_02162_),
    .A2(_02165_),
    .A3(_02168_),
    .B1(_09562_),
    .X(_02177_));
 sky130_fd_sc_hd__o211ai_2 _26327_ (.A1(_09553_),
    .A2(_09556_),
    .B1(_02171_),
    .C1(_02173_),
    .Y(_02178_));
 sky130_fd_sc_hd__a31o_2 _26328_ (.A1(_09563_),
    .A2(_02171_),
    .A3(_02173_),
    .B1(_02175_),
    .X(_02179_));
 sky130_fd_sc_hd__o31a_1 _26329_ (.A1(_09562_),
    .A2(_02169_),
    .A3(_02172_),
    .B1(_02176_),
    .X(_02180_));
 sky130_fd_sc_hd__a2bb2oi_2 _26330_ (.A1_N(_05760_),
    .A2_N(_05762_),
    .B1(_02176_),
    .B2(_02178_),
    .Y(_02182_));
 sky130_fd_sc_hd__o211ai_4 _26331_ (.A1(_02161_),
    .A2(_09563_),
    .B1(_05768_),
    .C1(_02174_),
    .Y(_02183_));
 sky130_fd_sc_hd__o21ai_1 _26332_ (.A1(_02169_),
    .A2(_02177_),
    .B1(_05767_),
    .Y(_02184_));
 sky130_fd_sc_hd__o311a_1 _26333_ (.A1(_09562_),
    .A2(_02169_),
    .A3(_02172_),
    .B1(_02176_),
    .C1(_05767_),
    .X(_02185_));
 sky130_fd_sc_hd__o211ai_4 _26334_ (.A1(_02169_),
    .A2(_02177_),
    .B1(_02176_),
    .C1(_05767_),
    .Y(_02186_));
 sky130_fd_sc_hd__o21a_1 _26335_ (.A1(_02175_),
    .A2(_02184_),
    .B1(_02183_),
    .X(_02187_));
 sky130_fd_sc_hd__o21ai_1 _26336_ (.A1(_02175_),
    .A2(_02184_),
    .B1(_02183_),
    .Y(_02188_));
 sky130_fd_sc_hd__and4_1 _26337_ (.A(_00853_),
    .B(_00854_),
    .C(_01202_),
    .D(_01204_),
    .X(_02189_));
 sky130_fd_sc_hd__nand4_1 _26338_ (.A(_00853_),
    .B(_00854_),
    .C(_01202_),
    .D(_01204_),
    .Y(_02190_));
 sky130_fd_sc_hd__a211oi_2 _26339_ (.A1(_01519_),
    .A2(_01534_),
    .B1(_02190_),
    .C1(_01538_),
    .Y(_02191_));
 sky130_fd_sc_hd__nand3_1 _26340_ (.A(_01540_),
    .B(_01876_),
    .C(_02189_),
    .Y(_02193_));
 sky130_fd_sc_hd__a21oi_1 _26341_ (.A1(_02191_),
    .A2(_01876_),
    .B1(_01877_),
    .Y(_02194_));
 sky130_fd_sc_hd__o211ai_4 _26342_ (.A1(_01880_),
    .A2(_01874_),
    .B1(_01878_),
    .C1(_02193_),
    .Y(_02195_));
 sky130_fd_sc_hd__and4_1 _26343_ (.A(_02189_),
    .B(_01539_),
    .C(_01537_),
    .D(_00862_),
    .X(_02196_));
 sky130_fd_sc_hd__o211ai_4 _26344_ (.A1(_05507_),
    .A2(_01870_),
    .B1(_02191_),
    .C1(_00862_),
    .Y(_02197_));
 sky130_fd_sc_hd__nand2_1 _26345_ (.A(_01879_),
    .B(_02196_),
    .Y(_02198_));
 sky130_fd_sc_hd__a22oi_1 _26346_ (.A1(_01879_),
    .A2(_02196_),
    .B1(_01883_),
    .B2(_02194_),
    .Y(_02199_));
 sky130_fd_sc_hd__o21ai_2 _26347_ (.A1(_01874_),
    .A2(_02197_),
    .B1(_02195_),
    .Y(_02200_));
 sky130_fd_sc_hd__a21oi_2 _26348_ (.A1(_02183_),
    .A2(_02186_),
    .B1(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__and3_1 _26349_ (.A(_02183_),
    .B(_02186_),
    .C(_02200_),
    .X(_02202_));
 sky130_fd_sc_hd__o22ai_2 _26350_ (.A1(net142),
    .A2(_09573_),
    .B1(_02188_),
    .B2(_02199_),
    .Y(_02204_));
 sky130_fd_sc_hd__a22o_2 _26351_ (.A1(_09575_),
    .A2(_09577_),
    .B1(_02176_),
    .B2(_02178_),
    .X(_02205_));
 sky130_fd_sc_hd__inv_2 _26352_ (.A(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__o21ai_2 _26353_ (.A1(_02182_),
    .A2(_02185_),
    .B1(_02200_),
    .Y(_02207_));
 sky130_fd_sc_hd__o211ai_4 _26354_ (.A1(_01874_),
    .A2(_02197_),
    .B1(_02195_),
    .C1(_02186_),
    .Y(_02208_));
 sky130_fd_sc_hd__o2111ai_4 _26355_ (.A1(_05768_),
    .A2(_02179_),
    .B1(_02183_),
    .C1(_02195_),
    .D1(_02198_),
    .Y(_02209_));
 sky130_fd_sc_hd__o221ai_4 _26356_ (.A1(net142),
    .A2(_09573_),
    .B1(_02182_),
    .B2(_02208_),
    .C1(_02207_),
    .Y(_02210_));
 sky130_fd_sc_hd__o221a_1 _26357_ (.A1(_09579_),
    .A2(_02179_),
    .B1(_02201_),
    .B2(_02204_),
    .C1(_10479_),
    .X(_02211_));
 sky130_fd_sc_hd__a211o_1 _26358_ (.A1(_02205_),
    .A2(_02210_),
    .B1(net141),
    .C1(_10475_),
    .X(_02212_));
 sky130_fd_sc_hd__a311oi_4 _26359_ (.A1(_09579_),
    .A2(_02207_),
    .A3(_02209_),
    .B1(_02206_),
    .C1(_05508_),
    .Y(_02213_));
 sky130_fd_sc_hd__nand3_4 _26360_ (.A(_02210_),
    .B(_05507_),
    .C(_02205_),
    .Y(_02215_));
 sky130_fd_sc_hd__a2bb2oi_1 _26361_ (.A1_N(_05500_),
    .A2_N(_05503_),
    .B1(_02205_),
    .B2(_02210_),
    .Y(_02216_));
 sky130_fd_sc_hd__o221ai_4 _26362_ (.A1(_09579_),
    .A2(_02179_),
    .B1(_02201_),
    .B2(_02204_),
    .C1(net292),
    .Y(_02217_));
 sky130_fd_sc_hd__o221a_1 _26363_ (.A1(_01555_),
    .A2(_01552_),
    .B1(_05248_),
    .B2(_01887_),
    .C1(_01550_),
    .X(_02218_));
 sky130_fd_sc_hd__a21oi_2 _26364_ (.A1(_01890_),
    .A2(_01892_),
    .B1(_01893_),
    .Y(_02219_));
 sky130_fd_sc_hd__o2bb2ai_1 _26365_ (.A1_N(_02215_),
    .A2_N(_02217_),
    .B1(_02218_),
    .B2(_01891_),
    .Y(_02220_));
 sky130_fd_sc_hd__nand3b_1 _26366_ (.A_N(_02219_),
    .B(_02217_),
    .C(_02215_),
    .Y(_02221_));
 sky130_fd_sc_hd__o311a_1 _26367_ (.A1(_02219_),
    .A2(_02216_),
    .A3(_02213_),
    .B1(net131),
    .C1(_02220_),
    .X(_02222_));
 sky130_fd_sc_hd__o211ai_2 _26368_ (.A1(net141),
    .A2(_10475_),
    .B1(_02220_),
    .C1(_02221_),
    .Y(_02223_));
 sky130_fd_sc_hd__a31o_2 _26369_ (.A1(net131),
    .A2(_02220_),
    .A3(_02221_),
    .B1(_02211_),
    .X(_02224_));
 sky130_fd_sc_hd__a2bb2oi_1 _26370_ (.A1_N(net318),
    .A2_N(net315),
    .B1(_02212_),
    .B2(_02223_),
    .Y(_02226_));
 sky130_fd_sc_hd__o22ai_2 _26371_ (.A1(net318),
    .A2(net315),
    .B1(_02211_),
    .B2(_02222_),
    .Y(_02227_));
 sky130_fd_sc_hd__o211a_1 _26372_ (.A1(_05246_),
    .A2(_05247_),
    .B1(_02212_),
    .C1(_02223_),
    .X(_02228_));
 sky130_fd_sc_hd__o211ai_2 _26373_ (.A1(_05246_),
    .A2(_05247_),
    .B1(_02212_),
    .C1(_02223_),
    .Y(_02229_));
 sky130_fd_sc_hd__o32a_1 _26374_ (.A1(net340),
    .A2(_04184_),
    .A3(_01900_),
    .B1(_01902_),
    .B2(_01598_),
    .X(_02230_));
 sky130_fd_sc_hd__o32ai_2 _26375_ (.A1(net340),
    .A2(_04184_),
    .A3(_01900_),
    .B1(_01902_),
    .B2(_01598_),
    .Y(_02231_));
 sky130_fd_sc_hd__nand3_1 _26376_ (.A(_02227_),
    .B(_02229_),
    .C(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__o21ai_1 _26377_ (.A1(_02226_),
    .A2(_02228_),
    .B1(_02230_),
    .Y(_02233_));
 sky130_fd_sc_hd__o211ai_2 _26378_ (.A1(net137),
    .A2(_10951_),
    .B1(_02232_),
    .C1(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__a211o_1 _26379_ (.A1(_02212_),
    .A2(_02223_),
    .B1(net137),
    .C1(_10951_),
    .X(_02235_));
 sky130_fd_sc_hd__o21ai_1 _26380_ (.A1(_02226_),
    .A2(_02228_),
    .B1(_02231_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand3_1 _26381_ (.A(_02230_),
    .B(_02229_),
    .C(_02227_),
    .Y(_02238_));
 sky130_fd_sc_hd__o211ai_1 _26382_ (.A1(net137),
    .A2(_10951_),
    .B1(_02237_),
    .C1(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__o21ai_1 _26383_ (.A1(_10954_),
    .A2(_02224_),
    .B1(_02234_),
    .Y(_02240_));
 sky130_fd_sc_hd__a31o_1 _26384_ (.A1(_01911_),
    .A2(_01914_),
    .A3(_01916_),
    .B1(_01907_),
    .X(_02241_));
 sky130_fd_sc_hd__a31oi_4 _26385_ (.A1(_01911_),
    .A2(_01914_),
    .A3(_01916_),
    .B1(_01907_),
    .Y(_02242_));
 sky130_fd_sc_hd__and3_1 _26386_ (.A(_02239_),
    .B(_04227_),
    .C(_02235_),
    .X(_02243_));
 sky130_fd_sc_hd__o211ai_2 _26387_ (.A1(_04206_),
    .A2(_04216_),
    .B1(_02235_),
    .C1(_02239_),
    .Y(_02244_));
 sky130_fd_sc_hd__o211ai_4 _26388_ (.A1(_10954_),
    .A2(_02224_),
    .B1(_02234_),
    .C1(_04238_),
    .Y(_02245_));
 sky130_fd_sc_hd__nand2_1 _26389_ (.A(_02244_),
    .B(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__nand3_1 _26390_ (.A(_02241_),
    .B(_02244_),
    .C(_02245_),
    .Y(_02248_));
 sky130_fd_sc_hd__nand2_1 _26391_ (.A(_02242_),
    .B(_02246_),
    .Y(_02249_));
 sky130_fd_sc_hd__o211ai_2 _26392_ (.A1(_11459_),
    .A2(_11461_),
    .B1(_02248_),
    .C1(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__o21ai_2 _26393_ (.A1(_11465_),
    .A2(_02240_),
    .B1(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__o21a_1 _26394_ (.A1(_02049_),
    .A2(net343),
    .B1(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__o311a_1 _26395_ (.A1(_11459_),
    .A2(net129),
    .A3(_02240_),
    .B1(_02137_),
    .C1(_02250_),
    .X(_02253_));
 sky130_fd_sc_hd__nor2_1 _26396_ (.A(_02252_),
    .B(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__a21oi_1 _26397_ (.A1(_01925_),
    .A2(_01926_),
    .B1(_01923_),
    .Y(_02255_));
 sky130_fd_sc_hd__a32o_1 _26398_ (.A1(_00240_),
    .A2(_01921_),
    .A3(_01922_),
    .B1(_01925_),
    .B2(_01926_),
    .X(_02256_));
 sky130_fd_sc_hd__o21ai_1 _26399_ (.A1(_02252_),
    .A2(_02253_),
    .B1(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__a21oi_1 _26400_ (.A1(_02257_),
    .A2(_11943_),
    .B1(_02251_),
    .Y(_02259_));
 sky130_fd_sc_hd__xnor2_1 _26401_ (.A(_01932_),
    .B(_02259_),
    .Y(net102));
 sky130_fd_sc_hd__a2111o_1 _26402_ (.A1(_11943_),
    .A2(_02257_),
    .B1(_02251_),
    .C1(_01928_),
    .D1(_01597_),
    .X(_02260_));
 sky130_fd_sc_hd__a31o_1 _26403_ (.A1(_01934_),
    .A2(_04029_),
    .A3(_10971_),
    .B1(_11470_),
    .X(_02261_));
 sky130_fd_sc_hd__o21ai_2 _26404_ (.A1(_02261_),
    .A2(_01942_),
    .B1(net271),
    .Y(_02262_));
 sky130_fd_sc_hd__o311a_1 _26405_ (.A1(_11470_),
    .A2(_01938_),
    .A3(_01942_),
    .B1(_05486_),
    .C1(net271),
    .X(_02263_));
 sky130_fd_sc_hd__or3_1 _26406_ (.A(net270),
    .B(net268),
    .C(_02262_),
    .X(_02264_));
 sky130_fd_sc_hd__o211ai_4 _26407_ (.A1(_02261_),
    .A2(_01942_),
    .B1(_10971_),
    .C1(net271),
    .Y(_02265_));
 sky130_fd_sc_hd__o21ai_2 _26408_ (.A1(_10965_),
    .A2(_10967_),
    .B1(_02262_),
    .Y(_02266_));
 sky130_fd_sc_hd__nand2_1 _26409_ (.A(_02265_),
    .B(_02266_),
    .Y(_02267_));
 sky130_fd_sc_hd__o221ai_4 _26410_ (.A1(net153),
    .A2(_01625_),
    .B1(_01946_),
    .B2(net150),
    .C1(_01952_),
    .Y(_02269_));
 sky130_fd_sc_hd__o2111ai_4 _26411_ (.A1(_01935_),
    .A2(_01949_),
    .B1(_02265_),
    .C1(_02266_),
    .D1(_02269_),
    .Y(_02270_));
 sky130_fd_sc_hd__o211ai_2 _26412_ (.A1(_01950_),
    .A2(_01954_),
    .B1(_02267_),
    .C1(_01948_),
    .Y(_02271_));
 sky130_fd_sc_hd__nand3_1 _26413_ (.A(_02271_),
    .B(net244),
    .C(_02270_),
    .Y(_02272_));
 sky130_fd_sc_hd__o21a_2 _26414_ (.A1(net244),
    .A2(_02262_),
    .B1(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__a31o_2 _26415_ (.A1(_02271_),
    .A2(net244),
    .A3(_02270_),
    .B1(_02263_),
    .X(_02274_));
 sky130_fd_sc_hd__a2bb2oi_1 _26416_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_02264_),
    .B2(_02272_),
    .Y(_02275_));
 sky130_fd_sc_hd__a2bb2o_1 _26417_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_02264_),
    .B2(_02272_),
    .X(_02276_));
 sky130_fd_sc_hd__a31oi_1 _26418_ (.A1(_02271_),
    .A2(net244),
    .A3(_02270_),
    .B1(_10492_),
    .Y(_02277_));
 sky130_fd_sc_hd__a31o_1 _26419_ (.A1(_02271_),
    .A2(net244),
    .A3(_02270_),
    .B1(_10492_),
    .X(_02278_));
 sky130_fd_sc_hd__and3_1 _26420_ (.A(_02272_),
    .B(net150),
    .C(_02264_),
    .X(_02280_));
 sky130_fd_sc_hd__a21oi_1 _26421_ (.A1(_02264_),
    .A2(_02277_),
    .B1(_02275_),
    .Y(_02281_));
 sky130_fd_sc_hd__o2bb2ai_1 _26422_ (.A1_N(_01974_),
    .A2_N(_01975_),
    .B1(net153),
    .B2(_01963_),
    .Y(_02282_));
 sky130_fd_sc_hd__o211ai_2 _26423_ (.A1(_01961_),
    .A2(net151),
    .B1(_01975_),
    .C1(_01974_),
    .Y(_02283_));
 sky130_fd_sc_hd__a31oi_4 _26424_ (.A1(_01967_),
    .A2(_01974_),
    .A3(_01975_),
    .B1(_01964_),
    .Y(_02284_));
 sky130_fd_sc_hd__o2111a_1 _26425_ (.A1(_02278_),
    .A2(_02263_),
    .B1(_01965_),
    .C1(_02276_),
    .D1(_02283_),
    .X(_02285_));
 sky130_fd_sc_hd__o22ai_2 _26426_ (.A1(net265),
    .A2(net264),
    .B1(_02281_),
    .B2(_02284_),
    .Y(_02286_));
 sky130_fd_sc_hd__o211ai_1 _26427_ (.A1(_02275_),
    .A2(_02280_),
    .B1(_01965_),
    .C1(_01979_),
    .Y(_02287_));
 sky130_fd_sc_hd__o211ai_1 _26428_ (.A1(net151),
    .A2(_01961_),
    .B1(_02281_),
    .C1(_02282_),
    .Y(_02288_));
 sky130_fd_sc_hd__or3_1 _26429_ (.A(net265),
    .B(net264),
    .C(_02273_),
    .X(_02289_));
 sky130_fd_sc_hd__nand3_2 _26430_ (.A(_02288_),
    .B(_05752_),
    .C(_02287_),
    .Y(_02291_));
 sky130_fd_sc_hd__o21ai_4 _26431_ (.A1(_05752_),
    .A2(_02273_),
    .B1(_02291_),
    .Y(_02292_));
 sky130_fd_sc_hd__inv_2 _26432_ (.A(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__o221ai_4 _26433_ (.A1(_05752_),
    .A2(_02274_),
    .B1(_02285_),
    .B2(_02286_),
    .C1(net151),
    .Y(_02294_));
 sky130_fd_sc_hd__nand3_1 _26434_ (.A(_02291_),
    .B(net153),
    .C(_02289_),
    .Y(_02295_));
 sky130_fd_sc_hd__nand2_1 _26435_ (.A(_02294_),
    .B(_02295_),
    .Y(_02296_));
 sky130_fd_sc_hd__and3_1 _26436_ (.A(_01354_),
    .B(_01355_),
    .C(_01016_),
    .X(_02297_));
 sky130_fd_sc_hd__nand4_1 _26437_ (.A(_01013_),
    .B(_01015_),
    .C(_01354_),
    .D(_01355_),
    .Y(_02298_));
 sky130_fd_sc_hd__a211oi_2 _26438_ (.A1(_01652_),
    .A2(_01672_),
    .B1(_02298_),
    .C1(_01675_),
    .Y(_02299_));
 sky130_fd_sc_hd__nand3_1 _26439_ (.A(_01988_),
    .B(_02297_),
    .C(_01678_),
    .Y(_02300_));
 sky130_fd_sc_hd__o211a_1 _26440_ (.A1(_01993_),
    .A2(_01987_),
    .B1(_01989_),
    .C1(_02300_),
    .X(_02302_));
 sky130_fd_sc_hd__o211ai_4 _26441_ (.A1(_01993_),
    .A2(_01987_),
    .B1(_01989_),
    .C1(_02300_),
    .Y(_02303_));
 sky130_fd_sc_hd__o211ai_2 _26442_ (.A1(_01023_),
    .A2(_01027_),
    .B1(_02299_),
    .C1(_01989_),
    .Y(_02304_));
 sky130_fd_sc_hd__nand4_4 _26443_ (.A(_02299_),
    .B(_01989_),
    .C(_01988_),
    .D(_01029_),
    .Y(_02305_));
 sky130_fd_sc_hd__a21oi_2 _26444_ (.A1(_02303_),
    .A2(_02305_),
    .B1(_02296_),
    .Y(_02306_));
 sky130_fd_sc_hd__a21o_1 _26445_ (.A1(_02303_),
    .A2(_02305_),
    .B1(_02296_),
    .X(_02307_));
 sky130_fd_sc_hd__o211ai_1 _26446_ (.A1(_02304_),
    .A2(_01987_),
    .B1(_02296_),
    .C1(_02303_),
    .Y(_02308_));
 sky130_fd_sc_hd__a31oi_1 _26447_ (.A1(_02296_),
    .A2(_02303_),
    .A3(_02305_),
    .B1(_05995_),
    .Y(_02309_));
 sky130_fd_sc_hd__o21ai_2 _26448_ (.A1(net260),
    .A2(net255),
    .B1(_02308_),
    .Y(_02310_));
 sky130_fd_sc_hd__o211ai_2 _26449_ (.A1(_01987_),
    .A2(_02304_),
    .B1(_02295_),
    .C1(_02294_),
    .Y(_02311_));
 sky130_fd_sc_hd__a22o_1 _26450_ (.A1(_02294_),
    .A2(_02295_),
    .B1(_02303_),
    .B2(_02305_),
    .X(_02313_));
 sky130_fd_sc_hd__a211o_1 _26451_ (.A1(_02289_),
    .A2(_02291_),
    .B1(net260),
    .C1(net255),
    .X(_02314_));
 sky130_fd_sc_hd__o221ai_4 _26452_ (.A1(net260),
    .A2(net255),
    .B1(_02302_),
    .B2(_02311_),
    .C1(_02313_),
    .Y(_02315_));
 sky130_fd_sc_hd__a2bb2oi_2 _26453_ (.A1_N(net240),
    .A2_N(_02292_),
    .B1(_02307_),
    .B2(_02309_),
    .Y(_02316_));
 sky130_fd_sc_hd__a22o_2 _26454_ (.A1(_05995_),
    .A2(_02293_),
    .B1(_02309_),
    .B2(_02307_),
    .X(_02317_));
 sky130_fd_sc_hd__o221a_1 _26455_ (.A1(net240),
    .A2(_02292_),
    .B1(_02306_),
    .B2(_02310_),
    .C1(_06294_),
    .X(_02318_));
 sky130_fd_sc_hd__inv_2 _26456_ (.A(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__nand3_4 _26457_ (.A(_02315_),
    .B(net172),
    .C(_02314_),
    .Y(_02320_));
 sky130_fd_sc_hd__o221ai_4 _26458_ (.A1(net240),
    .A2(_02292_),
    .B1(_02306_),
    .B2(_02310_),
    .C1(net171),
    .Y(_02321_));
 sky130_fd_sc_hd__o2bb2a_1 _26459_ (.A1_N(net173),
    .A2_N(_02000_),
    .B1(_02001_),
    .B2(_01691_),
    .X(_02322_));
 sky130_fd_sc_hd__o211a_1 _26460_ (.A1(net175),
    .A2(_01686_),
    .B1(_02002_),
    .C1(_02007_),
    .X(_02324_));
 sky130_fd_sc_hd__o211ai_1 _26461_ (.A1(_08731_),
    .A2(_01686_),
    .B1(_02002_),
    .C1(_02007_),
    .Y(_02325_));
 sky130_fd_sc_hd__o21ai_2 _26462_ (.A1(net174),
    .A2(_01999_),
    .B1(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__a21oi_4 _26463_ (.A1(_02320_),
    .A2(_02321_),
    .B1(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__o2bb2ai_1 _26464_ (.A1_N(_02320_),
    .A2_N(_02321_),
    .B1(_02322_),
    .B2(_02005_),
    .Y(_02328_));
 sky130_fd_sc_hd__o211a_1 _26465_ (.A1(_02008_),
    .A2(_02324_),
    .B1(_02321_),
    .C1(_02320_),
    .X(_02329_));
 sky130_fd_sc_hd__nand3_4 _26466_ (.A(_02320_),
    .B(_02326_),
    .C(_02321_),
    .Y(_02330_));
 sky130_fd_sc_hd__o21ai_2 _26467_ (.A1(net239),
    .A2(_06292_),
    .B1(_02330_),
    .Y(_02331_));
 sky130_fd_sc_hd__o211ai_1 _26468_ (.A1(net239),
    .A2(_06292_),
    .B1(_02328_),
    .C1(_02330_),
    .Y(_02332_));
 sky130_fd_sc_hd__o22ai_2 _26469_ (.A1(net239),
    .A2(_06292_),
    .B1(_02327_),
    .B2(_02329_),
    .Y(_02333_));
 sky130_fd_sc_hd__o22a_2 _26470_ (.A1(_06293_),
    .A2(_02317_),
    .B1(_02327_),
    .B2(_02331_),
    .X(_02335_));
 sky130_fd_sc_hd__a31o_1 _26471_ (.A1(_02328_),
    .A2(_02330_),
    .A3(_06293_),
    .B1(_02318_),
    .X(_02336_));
 sky130_fd_sc_hd__o221ai_4 _26472_ (.A1(net200),
    .A2(_01707_),
    .B1(_02022_),
    .B2(_01723_),
    .C1(_02017_),
    .Y(_02337_));
 sky130_fd_sc_hd__o21ai_1 _26473_ (.A1(_02018_),
    .A2(_02023_),
    .B1(_02017_),
    .Y(_02338_));
 sky130_fd_sc_hd__o21ai_1 _26474_ (.A1(_02327_),
    .A2(_02331_),
    .B1(_09139_),
    .Y(_02339_));
 sky130_fd_sc_hd__o221a_1 _26475_ (.A1(_06293_),
    .A2(_02317_),
    .B1(_02327_),
    .B2(_02331_),
    .C1(_09139_),
    .X(_02340_));
 sky130_fd_sc_hd__o221ai_4 _26476_ (.A1(_06293_),
    .A2(_02317_),
    .B1(_02327_),
    .B2(_02331_),
    .C1(_09139_),
    .Y(_02341_));
 sky130_fd_sc_hd__a2bb2oi_2 _26477_ (.A1_N(net194),
    .A2_N(net191),
    .B1(_02319_),
    .B2(_02332_),
    .Y(_02342_));
 sky130_fd_sc_hd__o221ai_4 _26478_ (.A1(net194),
    .A2(net192),
    .B1(_02316_),
    .B2(_06293_),
    .C1(_02333_),
    .Y(_02343_));
 sky130_fd_sc_hd__o2111ai_1 _26479_ (.A1(_02018_),
    .A2(_02023_),
    .B1(_02341_),
    .C1(_02343_),
    .D1(_02017_),
    .Y(_02344_));
 sky130_fd_sc_hd__o21ai_1 _26480_ (.A1(_02340_),
    .A2(_02342_),
    .B1(_02338_),
    .Y(_02346_));
 sky130_fd_sc_hd__o211ai_2 _26481_ (.A1(net238),
    .A2(net236),
    .B1(_02344_),
    .C1(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__nand4_2 _26482_ (.A(_02019_),
    .B(_02337_),
    .C(_02341_),
    .D(_02343_),
    .Y(_02348_));
 sky130_fd_sc_hd__o2bb2ai_1 _26483_ (.A1_N(_02019_),
    .A2_N(_02337_),
    .B1(_02340_),
    .B2(_02342_),
    .Y(_02349_));
 sky130_fd_sc_hd__o211ai_4 _26484_ (.A1(net238),
    .A2(net236),
    .B1(_02348_),
    .C1(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__o31a_2 _26485_ (.A1(net238),
    .A2(net236),
    .A3(_02335_),
    .B1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__o211ai_4 _26486_ (.A1(_02336_),
    .A2(net209),
    .B1(_08731_),
    .C1(_02347_),
    .Y(_02352_));
 sky130_fd_sc_hd__o211a_2 _26487_ (.A1(net209),
    .A2(_02335_),
    .B1(net178),
    .C1(_02350_),
    .X(_02353_));
 sky130_fd_sc_hd__o211ai_4 _26488_ (.A1(net209),
    .A2(_02335_),
    .B1(net178),
    .C1(_02350_),
    .Y(_02354_));
 sky130_fd_sc_hd__nand2_1 _26489_ (.A(_02352_),
    .B(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__o22a_1 _26490_ (.A1(_08314_),
    .A2(_02032_),
    .B1(_01739_),
    .B2(_02045_),
    .X(_02357_));
 sky130_fd_sc_hd__o211ai_2 _26491_ (.A1(_02045_),
    .A2(_01739_),
    .B1(_02036_),
    .C1(_02043_),
    .Y(_02358_));
 sky130_fd_sc_hd__a31oi_2 _26492_ (.A1(_02036_),
    .A2(_02043_),
    .A3(_02046_),
    .B1(_02033_),
    .Y(_02359_));
 sky130_fd_sc_hd__a221oi_4 _26493_ (.A1(_02357_),
    .A2(_02043_),
    .B1(_02352_),
    .B2(_02354_),
    .C1(_02033_),
    .Y(_02360_));
 sky130_fd_sc_hd__o22ai_4 _26494_ (.A1(net229),
    .A2(net228),
    .B1(_02355_),
    .B2(_02359_),
    .Y(_02361_));
 sky130_fd_sc_hd__o32a_2 _26495_ (.A1(net229),
    .A2(net228),
    .A3(_02351_),
    .B1(_02360_),
    .B2(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__o22ai_4 _26496_ (.A1(_06903_),
    .A2(_02351_),
    .B1(_02360_),
    .B2(_02361_),
    .Y(_02363_));
 sky130_fd_sc_hd__or3_2 _26497_ (.A(net207),
    .B(net204),
    .C(_02362_),
    .X(_02364_));
 sky130_fd_sc_hd__inv_2 _26498_ (.A(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__o21a_1 _26499_ (.A1(_08307_),
    .A2(net216),
    .B1(_02363_),
    .X(_02366_));
 sky130_fd_sc_hd__o21ai_2 _26500_ (.A1(_08307_),
    .A2(net216),
    .B1(_02363_),
    .Y(_02368_));
 sky130_fd_sc_hd__o221ai_4 _26501_ (.A1(_06903_),
    .A2(_02351_),
    .B1(_02360_),
    .B2(_02361_),
    .C1(net200),
    .Y(_02369_));
 sky130_fd_sc_hd__nand4_1 _26502_ (.A(_01082_),
    .B(_01083_),
    .C(_01426_),
    .D(_01428_),
    .Y(_02370_));
 sky130_fd_sc_hd__a211oi_2 _26503_ (.A1(_01738_),
    .A2(_01751_),
    .B1(_02370_),
    .C1(_01755_),
    .Y(_02371_));
 sky130_fd_sc_hd__nand2_1 _26504_ (.A(_02062_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__o211ai_4 _26505_ (.A1(_02066_),
    .A2(_02061_),
    .B1(_02063_),
    .C1(_02372_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand4_4 _26506_ (.A(_02371_),
    .B(_02063_),
    .C(_02062_),
    .D(_01091_),
    .Y(_02374_));
 sky130_fd_sc_hd__nand2_1 _26507_ (.A(_02373_),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__a22oi_2 _26508_ (.A1(_02368_),
    .A2(_02369_),
    .B1(_02373_),
    .B2(_02374_),
    .Y(_02376_));
 sky130_fd_sc_hd__a22o_1 _26509_ (.A1(_02368_),
    .A2(_02369_),
    .B1(_02373_),
    .B2(_02374_),
    .X(_02377_));
 sky130_fd_sc_hd__nand3_4 _26510_ (.A(_02369_),
    .B(_02373_),
    .C(_02374_),
    .Y(_02379_));
 sky130_fd_sc_hd__o2111a_1 _26511_ (.A1(_08314_),
    .A2(_02363_),
    .B1(_02368_),
    .C1(_02373_),
    .D1(_02374_),
    .X(_02380_));
 sky130_fd_sc_hd__nor3_2 _26512_ (.A(_07232_),
    .B(_02376_),
    .C(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__o221ai_4 _26513_ (.A1(net207),
    .A2(net205),
    .B1(_02366_),
    .B2(_02379_),
    .C1(_02377_),
    .Y(_02382_));
 sky130_fd_sc_hd__o211a_4 _26514_ (.A1(_02365_),
    .A2(_02381_),
    .B1(_07545_),
    .C1(_07547_),
    .X(_02383_));
 sky130_fd_sc_hd__a211o_2 _26515_ (.A1(_02364_),
    .A2(_02382_),
    .B1(_07544_),
    .C1(_07546_),
    .X(_02384_));
 sky130_fd_sc_hd__o311a_2 _26516_ (.A1(_07232_),
    .A2(_02376_),
    .A3(_02380_),
    .B1(_07935_),
    .C1(_02364_),
    .X(_02385_));
 sky130_fd_sc_hd__o211ai_4 _26517_ (.A1(_07233_),
    .A2(_02362_),
    .B1(_07935_),
    .C1(_02382_),
    .Y(_02386_));
 sky130_fd_sc_hd__a22oi_4 _26518_ (.A1(_07929_),
    .A2(_07932_),
    .B1(_02364_),
    .B2(_02382_),
    .Y(_02387_));
 sky130_fd_sc_hd__o22ai_4 _26519_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_02365_),
    .B2(_02381_),
    .Y(_02388_));
 sky130_fd_sc_hd__a31o_1 _26520_ (.A1(_01770_),
    .A2(_02076_),
    .A3(_02080_),
    .B1(_02081_),
    .X(_02390_));
 sky130_fd_sc_hd__a31oi_4 _26521_ (.A1(_01770_),
    .A2(_02076_),
    .A3(_02080_),
    .B1(_02081_),
    .Y(_02391_));
 sky130_fd_sc_hd__o21bai_4 _26522_ (.A1(_02385_),
    .A2(_02387_),
    .B1_N(_02390_),
    .Y(_02392_));
 sky130_fd_sc_hd__nand3_4 _26523_ (.A(_02386_),
    .B(_02388_),
    .C(_02390_),
    .Y(_02393_));
 sky130_fd_sc_hd__o311a_1 _26524_ (.A1(_02385_),
    .A2(_02387_),
    .A3(_02391_),
    .B1(_07548_),
    .C1(_02392_),
    .X(_02394_));
 sky130_fd_sc_hd__nand3_2 _26525_ (.A(_02392_),
    .B(_02393_),
    .C(_07548_),
    .Y(_02395_));
 sky130_fd_sc_hd__a31o_1 _26526_ (.A1(_02392_),
    .A2(_02393_),
    .A3(_07548_),
    .B1(_02383_),
    .X(_02396_));
 sky130_fd_sc_hd__o221a_1 _26527_ (.A1(_06922_),
    .A2(_01781_),
    .B1(_02091_),
    .B2(_07246_),
    .C1(_01803_),
    .X(_02397_));
 sky130_fd_sc_hd__o221ai_2 _26528_ (.A1(_06922_),
    .A2(_01781_),
    .B1(_07246_),
    .B2(_02091_),
    .C1(_01803_),
    .Y(_02398_));
 sky130_fd_sc_hd__a31oi_4 _26529_ (.A1(_01784_),
    .A2(_01803_),
    .A3(_02092_),
    .B1(_02094_),
    .Y(_02399_));
 sky130_fd_sc_hd__a31oi_1 _26530_ (.A1(_02392_),
    .A2(_02393_),
    .A3(_07548_),
    .B1(_07565_),
    .Y(_02401_));
 sky130_fd_sc_hd__a31o_1 _26531_ (.A1(_02392_),
    .A2(_02393_),
    .A3(_07548_),
    .B1(_07565_),
    .X(_02402_));
 sky130_fd_sc_hd__a311oi_4 _26532_ (.A1(_02392_),
    .A2(_02393_),
    .A3(_07548_),
    .B1(_07565_),
    .C1(_02383_),
    .Y(_02403_));
 sky130_fd_sc_hd__nand3_1 _26533_ (.A(_02395_),
    .B(_07564_),
    .C(_02384_),
    .Y(_02404_));
 sky130_fd_sc_hd__a2bb2oi_4 _26534_ (.A1_N(net221),
    .A2_N(net219),
    .B1(_02384_),
    .B2(_02395_),
    .Y(_02405_));
 sky130_fd_sc_hd__o22ai_4 _26535_ (.A1(net221),
    .A2(net220),
    .B1(_02383_),
    .B2(_02394_),
    .Y(_02406_));
 sky130_fd_sc_hd__a21oi_1 _26536_ (.A1(_02384_),
    .A2(_02401_),
    .B1(_02405_),
    .Y(_02407_));
 sky130_fd_sc_hd__o211ai_1 _26537_ (.A1(_02094_),
    .A2(_02397_),
    .B1(_02404_),
    .C1(_02406_),
    .Y(_02408_));
 sky130_fd_sc_hd__o21ai_1 _26538_ (.A1(_02403_),
    .A2(_02405_),
    .B1(_02399_),
    .Y(_02409_));
 sky130_fd_sc_hd__o211ai_2 _26539_ (.A1(net183),
    .A2(net182),
    .B1(_02408_),
    .C1(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__and3_1 _26540_ (.A(_07913_),
    .B(_07915_),
    .C(_02396_),
    .X(_02412_));
 sky130_fd_sc_hd__a211o_1 _26541_ (.A1(_02384_),
    .A2(_02395_),
    .B1(net183),
    .C1(net182),
    .X(_02413_));
 sky130_fd_sc_hd__o211ai_4 _26542_ (.A1(_02383_),
    .A2(_02402_),
    .B1(_02399_),
    .C1(_02406_),
    .Y(_02414_));
 sky130_fd_sc_hd__o22ai_4 _26543_ (.A1(_02094_),
    .A2(_02397_),
    .B1(_02403_),
    .B2(_02405_),
    .Y(_02415_));
 sky130_fd_sc_hd__o211ai_2 _26544_ (.A1(net183),
    .A2(net182),
    .B1(_02414_),
    .C1(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__a31oi_4 _26545_ (.A1(_02414_),
    .A2(_02415_),
    .A3(net162),
    .B1(_02412_),
    .Y(_02417_));
 sky130_fd_sc_hd__o211ai_4 _26546_ (.A1(_02396_),
    .A2(net162),
    .B1(net223),
    .C1(_02410_),
    .Y(_02418_));
 sky130_fd_sc_hd__and3_1 _26547_ (.A(_02416_),
    .B(_07246_),
    .C(_02413_),
    .X(_02419_));
 sky130_fd_sc_hd__o211ai_4 _26548_ (.A1(_07244_),
    .A2(net247),
    .B1(_02413_),
    .C1(_02416_),
    .Y(_02420_));
 sky130_fd_sc_hd__nand2_1 _26549_ (.A(_02418_),
    .B(_02420_),
    .Y(_02421_));
 sky130_fd_sc_hd__o22ai_1 _26550_ (.A1(_06922_),
    .A2(_02101_),
    .B1(_02120_),
    .B2(_02111_),
    .Y(_02423_));
 sky130_fd_sc_hd__a31oi_4 _26551_ (.A1(_02107_),
    .A2(_02112_),
    .A3(_02114_),
    .B1(_02105_),
    .Y(_02424_));
 sky130_fd_sc_hd__a221oi_4 _26552_ (.A1(_02119_),
    .A2(_02112_),
    .B1(_02420_),
    .B2(_02418_),
    .C1(_02105_),
    .Y(_02425_));
 sky130_fd_sc_hd__o221ai_2 _26553_ (.A1(_06922_),
    .A2(_02101_),
    .B1(_02111_),
    .B2(_02120_),
    .C1(_02421_),
    .Y(_02426_));
 sky130_fd_sc_hd__nand3_1 _26554_ (.A(_02423_),
    .B(_02420_),
    .C(_02418_),
    .Y(_02427_));
 sky130_fd_sc_hd__o22ai_4 _26555_ (.A1(net181),
    .A2(net179),
    .B1(_02421_),
    .B2(_02424_),
    .Y(_02428_));
 sky130_fd_sc_hd__o211ai_1 _26556_ (.A1(net181),
    .A2(net179),
    .B1(_02426_),
    .C1(_02427_),
    .Y(_02429_));
 sky130_fd_sc_hd__or3_2 _26557_ (.A(net181),
    .B(net179),
    .C(_02417_),
    .X(_02430_));
 sky130_fd_sc_hd__inv_2 _26558_ (.A(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__o32a_4 _26559_ (.A1(net181),
    .A2(net179),
    .A3(_02417_),
    .B1(_02425_),
    .B2(_02428_),
    .X(_02432_));
 sky130_fd_sc_hd__o21ai_4 _26560_ (.A1(_02425_),
    .A2(_02428_),
    .B1(_02430_),
    .Y(_02434_));
 sky130_fd_sc_hd__or3_2 _26561_ (.A(net157),
    .B(_08712_),
    .C(_02432_),
    .X(_02435_));
 sky130_fd_sc_hd__a22oi_2 _26562_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_02429_),
    .B2(_02430_),
    .Y(_02436_));
 sky130_fd_sc_hd__o21ai_4 _26563_ (.A1(_06914_),
    .A2(net250),
    .B1(_02434_),
    .Y(_02437_));
 sky130_fd_sc_hd__o22a_1 _26564_ (.A1(_06918_),
    .A2(net249),
    .B1(_02425_),
    .B2(_02428_),
    .X(_02438_));
 sky130_fd_sc_hd__a31o_2 _26565_ (.A1(_02427_),
    .A2(net159),
    .A3(_02426_),
    .B1(net226),
    .X(_02439_));
 sky130_fd_sc_hd__o221a_1 _26566_ (.A1(net159),
    .A2(_02417_),
    .B1(_02425_),
    .B2(_02428_),
    .C1(_06922_),
    .X(_02440_));
 sky130_fd_sc_hd__o221ai_4 _26567_ (.A1(net159),
    .A2(_02417_),
    .B1(_02425_),
    .B2(_02428_),
    .C1(_06922_),
    .Y(_02441_));
 sky130_fd_sc_hd__a21oi_1 _26568_ (.A1(_02430_),
    .A2(_02438_),
    .B1(_02436_),
    .Y(_02442_));
 sky130_fd_sc_hd__nand4_1 _26569_ (.A(_01159_),
    .B(_01161_),
    .C(_01489_),
    .D(_01490_),
    .Y(_02443_));
 sky130_fd_sc_hd__a211oi_1 _26570_ (.A1(_01807_),
    .A2(_01824_),
    .B1(_02443_),
    .C1(_01827_),
    .Y(_02445_));
 sky130_fd_sc_hd__nand2_1 _26571_ (.A(_02131_),
    .B(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__o211ai_4 _26572_ (.A1(_02135_),
    .A2(_02130_),
    .B1(_02133_),
    .C1(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__and4b_1 _26573_ (.A_N(_02443_),
    .B(_01828_),
    .C(_01826_),
    .D(_01164_),
    .X(_02448_));
 sky130_fd_sc_hd__o211ai_1 _26574_ (.A1(net235),
    .A2(_02125_),
    .B1(_02445_),
    .C1(_01164_),
    .Y(_02449_));
 sky130_fd_sc_hd__nand3_4 _26575_ (.A(_02448_),
    .B(_02133_),
    .C(_02131_),
    .Y(_02450_));
 sky130_fd_sc_hd__o21ai_2 _26576_ (.A1(_02130_),
    .A2(_02449_),
    .B1(_02447_),
    .Y(_02451_));
 sky130_fd_sc_hd__o211ai_1 _26577_ (.A1(_02436_),
    .A2(_02440_),
    .B1(_02447_),
    .C1(_02450_),
    .Y(_02452_));
 sky130_fd_sc_hd__nand2_1 _26578_ (.A(_02451_),
    .B(_02442_),
    .Y(_02453_));
 sky130_fd_sc_hd__a22o_1 _26579_ (.A1(_02437_),
    .A2(_02441_),
    .B1(_02447_),
    .B2(_02450_),
    .X(_02454_));
 sky130_fd_sc_hd__o2111ai_4 _26580_ (.A1(_02439_),
    .A2(_02431_),
    .B1(_02437_),
    .C1(_02447_),
    .D1(_02450_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand3_2 _26581_ (.A(_02454_),
    .B(_02456_),
    .C(net149),
    .Y(_02457_));
 sky130_fd_sc_hd__o221a_1 _26582_ (.A1(net159),
    .A2(_02417_),
    .B1(_02425_),
    .B2(_02428_),
    .C1(_08715_),
    .X(_02458_));
 sky130_fd_sc_hd__nand3_1 _26583_ (.A(_02453_),
    .B(net149),
    .C(_02452_),
    .Y(_02459_));
 sky130_fd_sc_hd__o21ai_4 _26584_ (.A1(net149),
    .A2(_02432_),
    .B1(_02457_),
    .Y(_02460_));
 sky130_fd_sc_hd__inv_2 _26585_ (.A(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__a311o_1 _26586_ (.A1(_02453_),
    .A2(net149),
    .A3(_02452_),
    .B1(_02458_),
    .C1(net146),
    .X(_02462_));
 sky130_fd_sc_hd__a31oi_2 _26587_ (.A1(_02454_),
    .A2(_02456_),
    .A3(net149),
    .B1(net233),
    .Y(_02463_));
 sky130_fd_sc_hd__nand3_4 _26588_ (.A(_02457_),
    .B(net235),
    .C(_02435_),
    .Y(_02464_));
 sky130_fd_sc_hd__inv_2 _26589_ (.A(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__o211ai_4 _26590_ (.A1(_02434_),
    .A2(net149),
    .B1(net233),
    .C1(_02459_),
    .Y(_02467_));
 sky130_fd_sc_hd__o2bb2a_1 _26591_ (.A1_N(net252),
    .A2_N(_02143_),
    .B1(_02144_),
    .B2(_01840_),
    .X(_02468_));
 sky130_fd_sc_hd__o21ai_2 _26592_ (.A1(_02146_),
    .A2(_02147_),
    .B1(_02151_),
    .Y(_02469_));
 sky130_fd_sc_hd__a21oi_2 _26593_ (.A1(_02149_),
    .A2(_02145_),
    .B1(_02150_),
    .Y(_02470_));
 sky130_fd_sc_hd__a21oi_1 _26594_ (.A1(_02464_),
    .A2(_02467_),
    .B1(_02469_),
    .Y(_02471_));
 sky130_fd_sc_hd__o2bb2ai_2 _26595_ (.A1_N(_02464_),
    .A2_N(_02467_),
    .B1(_02468_),
    .B2(_02147_),
    .Y(_02472_));
 sky130_fd_sc_hd__nand3_1 _26596_ (.A(_02464_),
    .B(_02467_),
    .C(_02469_),
    .Y(_02473_));
 sky130_fd_sc_hd__a31oi_2 _26597_ (.A1(_02464_),
    .A2(_02467_),
    .A3(_02469_),
    .B1(_09124_),
    .Y(_02474_));
 sky130_fd_sc_hd__a31o_1 _26598_ (.A1(_02464_),
    .A2(_02467_),
    .A3(_02469_),
    .B1(_09124_),
    .X(_02475_));
 sky130_fd_sc_hd__o211ai_2 _26599_ (.A1(net148),
    .A2(net147),
    .B1(_02472_),
    .C1(_02473_),
    .Y(_02476_));
 sky130_fd_sc_hd__o22ai_4 _26600_ (.A1(net146),
    .A2(_02461_),
    .B1(_02471_),
    .B2(_02475_),
    .Y(_02478_));
 sky130_fd_sc_hd__a21oi_1 _26601_ (.A1(_02161_),
    .A2(_06014_),
    .B1(_02168_),
    .Y(_02479_));
 sky130_fd_sc_hd__a31o_1 _26602_ (.A1(_06013_),
    .A2(_02156_),
    .A3(_02160_),
    .B1(_02167_),
    .X(_02480_));
 sky130_fd_sc_hd__a32oi_4 _26603_ (.A1(_06013_),
    .A2(_02156_),
    .A3(_02160_),
    .B1(_02162_),
    .B2(_02167_),
    .Y(_02481_));
 sky130_fd_sc_hd__o2bb2ai_1 _26604_ (.A1_N(_02167_),
    .A2_N(_02162_),
    .B1(_02155_),
    .B2(_02163_),
    .Y(_02482_));
 sky130_fd_sc_hd__a221oi_4 _26605_ (.A1(_09124_),
    .A2(_02460_),
    .B1(_02474_),
    .B2(_02472_),
    .C1(_06315_),
    .Y(_02483_));
 sky130_fd_sc_hd__nand3_1 _26606_ (.A(_02476_),
    .B(_06314_),
    .C(_02462_),
    .Y(_02484_));
 sky130_fd_sc_hd__a2bb2oi_2 _26607_ (.A1_N(net284),
    .A2_N(net281),
    .B1(_02462_),
    .B2(_02476_),
    .Y(_02485_));
 sky130_fd_sc_hd__o21ai_1 _26608_ (.A1(net284),
    .A2(net281),
    .B1(_02478_),
    .Y(_02486_));
 sky130_fd_sc_hd__o211ai_2 _26609_ (.A1(_02164_),
    .A2(_02479_),
    .B1(_02484_),
    .C1(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__o2bb2ai_1 _26610_ (.A1_N(_02162_),
    .A2_N(_02480_),
    .B1(_02483_),
    .B2(_02485_),
    .Y(_02489_));
 sky130_fd_sc_hd__o211ai_4 _26611_ (.A1(net156),
    .A2(_09556_),
    .B1(_02487_),
    .C1(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__a211o_1 _26612_ (.A1(_02462_),
    .A2(_02476_),
    .B1(net156),
    .C1(_09556_),
    .X(_02491_));
 sky130_fd_sc_hd__nand3_1 _26613_ (.A(_02486_),
    .B(_02481_),
    .C(_02484_),
    .Y(_02492_));
 sky130_fd_sc_hd__o22ai_2 _26614_ (.A1(_02164_),
    .A2(_02479_),
    .B1(_02483_),
    .B2(_02485_),
    .Y(_02493_));
 sky130_fd_sc_hd__o211ai_2 _26615_ (.A1(net156),
    .A2(_09556_),
    .B1(_02492_),
    .C1(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__nand2_1 _26616_ (.A(_02491_),
    .B(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__o21ai_4 _26617_ (.A1(_09563_),
    .A2(_02478_),
    .B1(_02490_),
    .Y(_02496_));
 sky130_fd_sc_hd__a2bb2oi_1 _26618_ (.A1_N(_06009_),
    .A2_N(net287),
    .B1(_02491_),
    .B2(_02494_),
    .Y(_02497_));
 sky130_fd_sc_hd__o211ai_4 _26619_ (.A1(_09563_),
    .A2(_02478_),
    .B1(_02490_),
    .C1(_06014_),
    .Y(_02498_));
 sky130_fd_sc_hd__a31oi_1 _26620_ (.A1(_09563_),
    .A2(_02492_),
    .A3(_02493_),
    .B1(_06014_),
    .Y(_02500_));
 sky130_fd_sc_hd__o211ai_2 _26621_ (.A1(net285),
    .A2(_06012_),
    .B1(_02491_),
    .C1(_02494_),
    .Y(_02501_));
 sky130_fd_sc_hd__a21oi_1 _26622_ (.A1(_02491_),
    .A2(_02500_),
    .B1(_02497_),
    .Y(_02502_));
 sky130_fd_sc_hd__a22oi_2 _26623_ (.A1(_02183_),
    .A2(_02208_),
    .B1(_02498_),
    .B2(_02501_),
    .Y(_02503_));
 sky130_fd_sc_hd__o2111a_1 _26624_ (.A1(_05767_),
    .A2(_02180_),
    .B1(_02208_),
    .C1(_02498_),
    .D1(_02501_),
    .X(_02504_));
 sky130_fd_sc_hd__o21ai_4 _26625_ (.A1(_02503_),
    .A2(_02504_),
    .B1(net132),
    .Y(_02505_));
 sky130_fd_sc_hd__or3_2 _26626_ (.A(net142),
    .B(_09573_),
    .C(_02496_),
    .X(_02506_));
 sky130_fd_sc_hd__o31a_2 _26627_ (.A1(net142),
    .A2(_09573_),
    .A3(_02496_),
    .B1(_02505_),
    .X(_02507_));
 sky130_fd_sc_hd__a21oi_2 _26628_ (.A1(_02505_),
    .A2(_02506_),
    .B1(net131),
    .Y(_02508_));
 sky130_fd_sc_hd__or3_1 _26629_ (.A(net141),
    .B(_10475_),
    .C(_02507_),
    .X(_02509_));
 sky130_fd_sc_hd__a21oi_4 _26630_ (.A1(_02505_),
    .A2(_02506_),
    .B1(_05767_),
    .Y(_02511_));
 sky130_fd_sc_hd__a22o_1 _26631_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_02505_),
    .B2(_02506_),
    .X(_02512_));
 sky130_fd_sc_hd__o221a_1 _26632_ (.A1(_05765_),
    .A2(net288),
    .B1(net132),
    .B2(_02496_),
    .C1(_02505_),
    .X(_02513_));
 sky130_fd_sc_hd__o221ai_4 _26633_ (.A1(_05765_),
    .A2(net288),
    .B1(net132),
    .B2(_02496_),
    .C1(_02505_),
    .Y(_02514_));
 sky130_fd_sc_hd__o2111ai_4 _26634_ (.A1(_01544_),
    .A2(_01551_),
    .B1(_01550_),
    .C1(_01214_),
    .D1(_01218_),
    .Y(_02515_));
 sky130_fd_sc_hd__a21oi_2 _26635_ (.A1(_05249_),
    .A2(_01888_),
    .B1(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__nor3_1 _26636_ (.A(_01891_),
    .B(_02515_),
    .C(_01893_),
    .Y(_02517_));
 sky130_fd_sc_hd__o211ai_2 _26637_ (.A1(_05249_),
    .A2(_01888_),
    .B1(_02516_),
    .C1(_02215_),
    .Y(_02518_));
 sky130_fd_sc_hd__o211ai_4 _26638_ (.A1(_02219_),
    .A2(_02213_),
    .B1(_02217_),
    .C1(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__o2111ai_4 _26639_ (.A1(_05249_),
    .A2(_01888_),
    .B1(_02215_),
    .C1(_02516_),
    .D1(_02217_),
    .Y(_02520_));
 sky130_fd_sc_hd__nand4_2 _26640_ (.A(_02517_),
    .B(_02217_),
    .C(_02215_),
    .D(_01226_),
    .Y(_02522_));
 sky130_fd_sc_hd__o21ai_4 _26641_ (.A1(_01227_),
    .A2(_02520_),
    .B1(_02519_),
    .Y(_02523_));
 sky130_fd_sc_hd__o21ai_4 _26642_ (.A1(_02511_),
    .A2(_02513_),
    .B1(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__o211ai_4 _26643_ (.A1(_01227_),
    .A2(_02520_),
    .B1(_02519_),
    .C1(_02514_),
    .Y(_02525_));
 sky130_fd_sc_hd__o2111ai_4 _26644_ (.A1(_01227_),
    .A2(_02520_),
    .B1(_02519_),
    .C1(_02514_),
    .D1(_02512_),
    .Y(_02526_));
 sky130_fd_sc_hd__o221a_1 _26645_ (.A1(net141),
    .A2(net140),
    .B1(_02511_),
    .B2(_02525_),
    .C1(_02524_),
    .X(_02527_));
 sky130_fd_sc_hd__o221ai_4 _26646_ (.A1(net141),
    .A2(_10475_),
    .B1(_02511_),
    .B2(_02525_),
    .C1(_02524_),
    .Y(_02528_));
 sky130_fd_sc_hd__a31oi_4 _26647_ (.A1(net131),
    .A2(_02524_),
    .A3(_02526_),
    .B1(_02508_),
    .Y(_02529_));
 sky130_fd_sc_hd__a21oi_1 _26648_ (.A1(_05249_),
    .A2(_02224_),
    .B1(_02230_),
    .Y(_02530_));
 sky130_fd_sc_hd__o32a_1 _26649_ (.A1(net318),
    .A2(net315),
    .A3(_02224_),
    .B1(_02226_),
    .B2(_02230_),
    .X(_02531_));
 sky130_fd_sc_hd__a21oi_1 _26650_ (.A1(_02230_),
    .A2(_02229_),
    .B1(_02226_),
    .Y(_02533_));
 sky130_fd_sc_hd__o311a_2 _26651_ (.A1(net141),
    .A2(_10475_),
    .A3(_02507_),
    .B1(_05507_),
    .C1(_02528_),
    .X(_02534_));
 sky130_fd_sc_hd__o2111ai_4 _26652_ (.A1(_02507_),
    .A2(net131),
    .B1(_05504_),
    .C1(_05502_),
    .D1(_02528_),
    .Y(_02535_));
 sky130_fd_sc_hd__a21oi_1 _26653_ (.A1(_02509_),
    .A2(_02528_),
    .B1(_05507_),
    .Y(_02536_));
 sky130_fd_sc_hd__o22ai_4 _26654_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_02508_),
    .B2(_02527_),
    .Y(_02537_));
 sky130_fd_sc_hd__o21ai_1 _26655_ (.A1(_05507_),
    .A2(_02529_),
    .B1(_02531_),
    .Y(_02538_));
 sky130_fd_sc_hd__o22ai_2 _26656_ (.A1(_02228_),
    .A2(_02530_),
    .B1(_02534_),
    .B2(_02536_),
    .Y(_02539_));
 sky130_fd_sc_hd__or3_1 _26657_ (.A(net137),
    .B(_10951_),
    .C(_02529_),
    .X(_02540_));
 sky130_fd_sc_hd__o221ai_4 _26658_ (.A1(net137),
    .A2(_10951_),
    .B1(_02534_),
    .B2(_02538_),
    .C1(_02539_),
    .Y(_02541_));
 sky130_fd_sc_hd__a21oi_1 _26659_ (.A1(_02540_),
    .A2(_02541_),
    .B1(_11465_),
    .Y(_02542_));
 sky130_fd_sc_hd__a2bb2oi_2 _26660_ (.A1_N(net318),
    .A2_N(net315),
    .B1(_02540_),
    .B2(_02541_),
    .Y(_02544_));
 sky130_fd_sc_hd__a22o_1 _26661_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_02540_),
    .B2(_02541_),
    .X(_02545_));
 sky130_fd_sc_hd__o211a_1 _26662_ (.A1(_10954_),
    .A2(_02529_),
    .B1(_05248_),
    .C1(_02541_),
    .X(_02546_));
 sky130_fd_sc_hd__o2111ai_4 _26663_ (.A1(_02529_),
    .A2(_10954_),
    .B1(_05245_),
    .C1(_05243_),
    .D1(_02541_),
    .Y(_02547_));
 sky130_fd_sc_hd__nor2_1 _26664_ (.A(_02544_),
    .B(_02546_),
    .Y(_02548_));
 sky130_fd_sc_hd__o21ai_2 _26665_ (.A1(_02243_),
    .A2(_02242_),
    .B1(_02245_),
    .Y(_02549_));
 sky130_fd_sc_hd__o221ai_2 _26666_ (.A1(_02242_),
    .A2(_02243_),
    .B1(_02544_),
    .B2(_02546_),
    .C1(_02245_),
    .Y(_02550_));
 sky130_fd_sc_hd__a31oi_2 _26667_ (.A1(_02545_),
    .A2(_02547_),
    .A3(_02549_),
    .B1(_11464_),
    .Y(_02551_));
 sky130_fd_sc_hd__a21o_1 _26668_ (.A1(_02551_),
    .A2(_02550_),
    .B1(_02542_),
    .X(_02552_));
 sky130_fd_sc_hd__a211oi_2 _26669_ (.A1(_02551_),
    .A2(_02550_),
    .B1(_02542_),
    .C1(_04238_),
    .Y(_02553_));
 sky130_fd_sc_hd__o21a_1 _26670_ (.A1(net340),
    .A2(_04184_),
    .B1(_02552_),
    .X(_02555_));
 sky130_fd_sc_hd__o21ai_1 _26671_ (.A1(net340),
    .A2(_04184_),
    .B1(_02552_),
    .Y(_02556_));
 sky130_fd_sc_hd__o32ai_4 _26672_ (.A1(_02049_),
    .A2(net343),
    .A3(_02251_),
    .B1(_02252_),
    .B2(_02255_),
    .Y(_02557_));
 sky130_fd_sc_hd__o21ai_1 _26673_ (.A1(_02553_),
    .A2(_02555_),
    .B1(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__a21o_1 _26674_ (.A1(_02558_),
    .A2(_11943_),
    .B1(_02552_),
    .X(_02559_));
 sky130_fd_sc_hd__a21oi_1 _26675_ (.A1(_05119_),
    .A2(_02260_),
    .B1(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__and3_1 _26676_ (.A(_05119_),
    .B(_02260_),
    .C(_02559_),
    .X(_02561_));
 sky130_fd_sc_hd__nor2_1 _26677_ (.A(_02560_),
    .B(_02561_),
    .Y(net103));
 sky130_fd_sc_hd__or4b_1 _26678_ (.A(_01597_),
    .B(_01928_),
    .C(_02559_),
    .D_N(_02259_),
    .X(_02562_));
 sky130_fd_sc_hd__o211ai_2 _26679_ (.A1(_02262_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_02270_),
    .Y(_02563_));
 sky130_fd_sc_hd__and3_1 _26680_ (.A(_02563_),
    .B(net244),
    .C(_05754_),
    .X(_02565_));
 sky130_fd_sc_hd__a311o_1 _26681_ (.A1(_11471_),
    .A2(_02265_),
    .A3(_02270_),
    .B1(_05752_),
    .C1(_05486_),
    .X(_02566_));
 sky130_fd_sc_hd__and3_2 _26682_ (.A(_02563_),
    .B(net244),
    .C(_10971_),
    .X(_02567_));
 sky130_fd_sc_hd__a311o_1 _26683_ (.A1(_11471_),
    .A2(_02265_),
    .A3(_02270_),
    .B1(_10970_),
    .C1(_05486_),
    .X(_02568_));
 sky130_fd_sc_hd__a21oi_2 _26684_ (.A1(_02563_),
    .A2(net244),
    .B1(_10971_),
    .Y(_02569_));
 sky130_fd_sc_hd__nor2_1 _26685_ (.A(_02567_),
    .B(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__o221ai_4 _26686_ (.A1(net153),
    .A2(_01963_),
    .B1(_02273_),
    .B2(net150),
    .C1(_02283_),
    .Y(_02571_));
 sky130_fd_sc_hd__o311a_1 _26687_ (.A1(_10487_),
    .A2(net166),
    .A3(_02274_),
    .B1(_02570_),
    .C1(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__o211ai_4 _26688_ (.A1(_10492_),
    .A2(_02274_),
    .B1(_02570_),
    .C1(_02571_),
    .Y(_02573_));
 sky130_fd_sc_hd__o221a_1 _26689_ (.A1(_02567_),
    .A2(_02569_),
    .B1(_02280_),
    .B2(_02284_),
    .C1(_02276_),
    .X(_02574_));
 sky130_fd_sc_hd__o221ai_4 _26690_ (.A1(_02567_),
    .A2(_02569_),
    .B1(_02280_),
    .B2(_02284_),
    .C1(_02276_),
    .Y(_02576_));
 sky130_fd_sc_hd__o211ai_1 _26691_ (.A1(net265),
    .A2(net264),
    .B1(_02573_),
    .C1(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__a211o_1 _26692_ (.A1(_02563_),
    .A2(net244),
    .B1(net265),
    .C1(net264),
    .X(_02578_));
 sky130_fd_sc_hd__o22ai_1 _26693_ (.A1(net265),
    .A2(net264),
    .B1(_02572_),
    .B2(_02574_),
    .Y(_02579_));
 sky130_fd_sc_hd__o31a_2 _26694_ (.A1(_05754_),
    .A2(_02572_),
    .A3(_02574_),
    .B1(_02566_),
    .X(_02580_));
 sky130_fd_sc_hd__a311o_1 _26695_ (.A1(_02576_),
    .A2(_05752_),
    .A3(_02573_),
    .B1(net240),
    .C1(_02565_),
    .X(_02581_));
 sky130_fd_sc_hd__a2bb2oi_2 _26696_ (.A1_N(_10487_),
    .A2_N(net166),
    .B1(_02566_),
    .B2(_02577_),
    .Y(_02582_));
 sky130_fd_sc_hd__o211ai_1 _26697_ (.A1(_10487_),
    .A2(net166),
    .B1(_02578_),
    .C1(_02579_),
    .Y(_02583_));
 sky130_fd_sc_hd__a31oi_1 _26698_ (.A1(_02576_),
    .A2(_05752_),
    .A3(_02573_),
    .B1(_10492_),
    .Y(_02584_));
 sky130_fd_sc_hd__a311o_1 _26699_ (.A1(_02576_),
    .A2(_05752_),
    .A3(_02573_),
    .B1(_10492_),
    .C1(_02565_),
    .X(_02585_));
 sky130_fd_sc_hd__a21oi_1 _26700_ (.A1(_02566_),
    .A2(_02584_),
    .B1(_02582_),
    .Y(_02587_));
 sky130_fd_sc_hd__nand2_1 _26701_ (.A(_02583_),
    .B(_02585_),
    .Y(_02588_));
 sky130_fd_sc_hd__o2bb2ai_1 _26702_ (.A1_N(_02303_),
    .A2_N(_02305_),
    .B1(net153),
    .B2(_02293_),
    .Y(_02589_));
 sky130_fd_sc_hd__o21ai_1 _26703_ (.A1(net151),
    .A2(_02292_),
    .B1(_02305_),
    .Y(_02590_));
 sky130_fd_sc_hd__o211ai_4 _26704_ (.A1(_02292_),
    .A2(net151),
    .B1(_02305_),
    .C1(_02303_),
    .Y(_02591_));
 sky130_fd_sc_hd__o22ai_2 _26705_ (.A1(net153),
    .A2(_02293_),
    .B1(_02590_),
    .B2(_02302_),
    .Y(_02592_));
 sky130_fd_sc_hd__o2111ai_1 _26706_ (.A1(net153),
    .A2(_02293_),
    .B1(_02583_),
    .C1(_02585_),
    .D1(_02591_),
    .Y(_02593_));
 sky130_fd_sc_hd__o211ai_1 _26707_ (.A1(net151),
    .A2(_02292_),
    .B1(_02588_),
    .C1(_02589_),
    .Y(_02594_));
 sky130_fd_sc_hd__a21oi_2 _26708_ (.A1(_02294_),
    .A2(_02591_),
    .B1(_02588_),
    .Y(_02595_));
 sky130_fd_sc_hd__o211ai_1 _26709_ (.A1(net260),
    .A2(net255),
    .B1(_02593_),
    .C1(_02594_),
    .Y(_02596_));
 sky130_fd_sc_hd__and3_1 _26710_ (.A(_02579_),
    .B(_05995_),
    .C(_02578_),
    .X(_02598_));
 sky130_fd_sc_hd__o22ai_4 _26711_ (.A1(net260),
    .A2(net255),
    .B1(_02587_),
    .B2(_02592_),
    .Y(_02599_));
 sky130_fd_sc_hd__o22ai_4 _26712_ (.A1(net240),
    .A2(_02580_),
    .B1(_02595_),
    .B2(_02599_),
    .Y(_02600_));
 sky130_fd_sc_hd__inv_2 _26713_ (.A(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__o21ai_4 _26714_ (.A1(_06286_),
    .A2(_06288_),
    .B1(_02600_),
    .Y(_02602_));
 sky130_fd_sc_hd__inv_2 _26715_ (.A(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__o211ai_2 _26716_ (.A1(net170),
    .A2(net168),
    .B1(_02581_),
    .C1(_02596_),
    .Y(_02604_));
 sky130_fd_sc_hd__o22ai_1 _26717_ (.A1(net167),
    .A2(_10024_),
    .B1(_02595_),
    .B2(_02599_),
    .Y(_02605_));
 sky130_fd_sc_hd__o21a_1 _26718_ (.A1(_02598_),
    .A2(_02605_),
    .B1(_02604_),
    .X(_02606_));
 sky130_fd_sc_hd__o21ai_1 _26719_ (.A1(_02598_),
    .A2(_02605_),
    .B1(_02604_),
    .Y(_02607_));
 sky130_fd_sc_hd__o2111ai_2 _26720_ (.A1(_01375_),
    .A2(_01366_),
    .B1(_01373_),
    .C1(_01690_),
    .D1(_01692_),
    .Y(_02609_));
 sky130_fd_sc_hd__a211oi_2 _26721_ (.A1(_01986_),
    .A2(_02004_),
    .B1(_02609_),
    .C1(_02008_),
    .Y(_02610_));
 sky130_fd_sc_hd__o21ai_2 _26722_ (.A1(net171),
    .A2(_02316_),
    .B1(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__o211a_1 _26723_ (.A1(_02317_),
    .A2(net172),
    .B1(_02611_),
    .C1(_02330_),
    .X(_02612_));
 sky130_fd_sc_hd__o211ai_4 _26724_ (.A1(_02317_),
    .A2(net172),
    .B1(_02611_),
    .C1(_02330_),
    .Y(_02613_));
 sky130_fd_sc_hd__nand4_4 _26725_ (.A(_02320_),
    .B(_02610_),
    .C(_02321_),
    .D(_01386_),
    .Y(_02614_));
 sky130_fd_sc_hd__nand3_1 _26726_ (.A(_02607_),
    .B(_02613_),
    .C(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__a21o_1 _26727_ (.A1(_02613_),
    .A2(_02614_),
    .B1(_02607_),
    .X(_02616_));
 sky130_fd_sc_hd__nand3_4 _26728_ (.A(_02606_),
    .B(_02613_),
    .C(_02614_),
    .Y(_02617_));
 sky130_fd_sc_hd__a21o_1 _26729_ (.A1(_02613_),
    .A2(_02614_),
    .B1(_02606_),
    .X(_02618_));
 sky130_fd_sc_hd__nand3_2 _26730_ (.A(_02618_),
    .B(_06293_),
    .C(_02617_),
    .Y(_02620_));
 sky130_fd_sc_hd__o221a_1 _26731_ (.A1(net240),
    .A2(_02580_),
    .B1(_02595_),
    .B2(_02599_),
    .C1(_06294_),
    .X(_02621_));
 sky130_fd_sc_hd__or3_1 _26732_ (.A(net239),
    .B(_06292_),
    .C(_02600_),
    .X(_02622_));
 sky130_fd_sc_hd__nand3_2 _26733_ (.A(_02616_),
    .B(_06293_),
    .C(_02615_),
    .Y(_02623_));
 sky130_fd_sc_hd__a31o_1 _26734_ (.A1(_02618_),
    .A2(_06293_),
    .A3(_02617_),
    .B1(_02603_),
    .X(_02624_));
 sky130_fd_sc_hd__o221a_4 _26735_ (.A1(_06605_),
    .A2(_06606_),
    .B1(_02600_),
    .B2(_06293_),
    .C1(_02623_),
    .X(_02625_));
 sky130_fd_sc_hd__a311o_2 _26736_ (.A1(_02616_),
    .A2(_06293_),
    .A3(_02615_),
    .B1(_02621_),
    .C1(net209),
    .X(_02626_));
 sky130_fd_sc_hd__a311oi_2 _26737_ (.A1(_02618_),
    .A2(_06293_),
    .A3(_02617_),
    .B1(net171),
    .C1(_02603_),
    .Y(_02627_));
 sky130_fd_sc_hd__nand3_4 _26738_ (.A(_02620_),
    .B(net172),
    .C(_02602_),
    .Y(_02628_));
 sky130_fd_sc_hd__a311oi_1 _26739_ (.A1(_02616_),
    .A2(_06293_),
    .A3(_02615_),
    .B1(_02621_),
    .C1(net172),
    .Y(_02629_));
 sky130_fd_sc_hd__o211ai_4 _26740_ (.A1(net189),
    .A2(net188),
    .B1(_02622_),
    .C1(_02623_),
    .Y(_02631_));
 sky130_fd_sc_hd__o221a_1 _26741_ (.A1(_02023_),
    .A2(_02018_),
    .B1(_09139_),
    .B2(_02335_),
    .C1(_02017_),
    .X(_02632_));
 sky130_fd_sc_hd__a22o_1 _26742_ (.A1(net173),
    .A2(_02336_),
    .B1(_02337_),
    .B2(_02019_),
    .X(_02633_));
 sky130_fd_sc_hd__a31o_1 _26743_ (.A1(_02019_),
    .A2(_02337_),
    .A3(_02341_),
    .B1(_02342_),
    .X(_02634_));
 sky130_fd_sc_hd__a31oi_2 _26744_ (.A1(_02019_),
    .A2(_02337_),
    .A3(_02341_),
    .B1(_02342_),
    .Y(_02635_));
 sky130_fd_sc_hd__a21oi_1 _26745_ (.A1(_02628_),
    .A2(_02631_),
    .B1(_02634_),
    .Y(_02636_));
 sky130_fd_sc_hd__o2bb2ai_4 _26746_ (.A1_N(_02628_),
    .A2_N(_02631_),
    .B1(_02632_),
    .B2(_02340_),
    .Y(_02637_));
 sky130_fd_sc_hd__o2111a_1 _26747_ (.A1(net173),
    .A2(_02336_),
    .B1(_02628_),
    .C1(_02631_),
    .D1(_02633_),
    .X(_02638_));
 sky130_fd_sc_hd__nand4_4 _26748_ (.A(_02341_),
    .B(_02628_),
    .C(_02631_),
    .D(_02633_),
    .Y(_02639_));
 sky130_fd_sc_hd__nand3_1 _26749_ (.A(_02637_),
    .B(_02639_),
    .C(net209),
    .Y(_02640_));
 sky130_fd_sc_hd__o22ai_2 _26750_ (.A1(net238),
    .A2(net236),
    .B1(_02636_),
    .B2(_02638_),
    .Y(_02642_));
 sky130_fd_sc_hd__o31a_1 _26751_ (.A1(_06613_),
    .A2(_02636_),
    .A3(_02638_),
    .B1(_02626_),
    .X(_02643_));
 sky130_fd_sc_hd__a31o_1 _26752_ (.A1(_02637_),
    .A2(_02639_),
    .A3(net209),
    .B1(_02625_),
    .X(_02644_));
 sky130_fd_sc_hd__o311a_1 _26753_ (.A1(_08311_),
    .A2(net215),
    .A3(_02031_),
    .B1(_02352_),
    .C1(_02358_),
    .X(_02645_));
 sky130_fd_sc_hd__a31oi_4 _26754_ (.A1(_02034_),
    .A2(_02352_),
    .A3(_02358_),
    .B1(_02353_),
    .Y(_02646_));
 sky130_fd_sc_hd__a31oi_1 _26755_ (.A1(_02637_),
    .A2(_02639_),
    .A3(net209),
    .B1(net173),
    .Y(_02647_));
 sky130_fd_sc_hd__a31o_2 _26756_ (.A1(_02637_),
    .A2(_02639_),
    .A3(net209),
    .B1(net173),
    .X(_02648_));
 sky130_fd_sc_hd__a311oi_4 _26757_ (.A1(_02637_),
    .A2(_02639_),
    .A3(net209),
    .B1(net173),
    .C1(_02625_),
    .Y(_02649_));
 sky130_fd_sc_hd__nand3_1 _26758_ (.A(_02640_),
    .B(_09139_),
    .C(_02626_),
    .Y(_02650_));
 sky130_fd_sc_hd__a2bb2oi_4 _26759_ (.A1_N(net194),
    .A2_N(net191),
    .B1(_02626_),
    .B2(_02640_),
    .Y(_02651_));
 sky130_fd_sc_hd__o221ai_4 _26760_ (.A1(net194),
    .A2(net191),
    .B1(_02624_),
    .B2(net209),
    .C1(_02642_),
    .Y(_02653_));
 sky130_fd_sc_hd__o221ai_2 _26761_ (.A1(_02353_),
    .A2(_02645_),
    .B1(_02648_),
    .B2(_02625_),
    .C1(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__o21ai_1 _26762_ (.A1(_02649_),
    .A2(_02651_),
    .B1(_02646_),
    .Y(_02655_));
 sky130_fd_sc_hd__o211ai_2 _26763_ (.A1(net229),
    .A2(net228),
    .B1(_02654_),
    .C1(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__o311a_1 _26764_ (.A1(net238),
    .A2(_02624_),
    .A3(net236),
    .B1(_06904_),
    .C1(_02642_),
    .X(_02657_));
 sky130_fd_sc_hd__o211ai_4 _26765_ (.A1(_02625_),
    .A2(_02648_),
    .B1(_02646_),
    .C1(_02653_),
    .Y(_02658_));
 sky130_fd_sc_hd__o22ai_4 _26766_ (.A1(_02353_),
    .A2(_02645_),
    .B1(_02649_),
    .B2(_02651_),
    .Y(_02659_));
 sky130_fd_sc_hd__o211ai_2 _26767_ (.A1(net229),
    .A2(net228),
    .B1(_02658_),
    .C1(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__a31oi_4 _26768_ (.A1(_02658_),
    .A2(_02659_),
    .A3(_06903_),
    .B1(_02657_),
    .Y(_02661_));
 sky130_fd_sc_hd__inv_2 _26769_ (.A(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__o211ai_4 _26770_ (.A1(_02644_),
    .A2(_06903_),
    .B1(_08731_),
    .C1(_02656_),
    .Y(_02664_));
 sky130_fd_sc_hd__o211a_1 _26771_ (.A1(_06903_),
    .A2(_02643_),
    .B1(net178),
    .C1(_02660_),
    .X(_02665_));
 sky130_fd_sc_hd__o211ai_2 _26772_ (.A1(_06903_),
    .A2(_02643_),
    .B1(net178),
    .C1(_02660_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_1 _26773_ (.A(_02664_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__a22o_1 _26774_ (.A1(_08314_),
    .A2(_02363_),
    .B1(_02373_),
    .B2(_02374_),
    .X(_02668_));
 sky130_fd_sc_hd__o2111ai_1 _26775_ (.A1(net200),
    .A2(_02362_),
    .B1(_02379_),
    .C1(_02664_),
    .D1(_02666_),
    .Y(_02669_));
 sky130_fd_sc_hd__o211ai_1 _26776_ (.A1(_08314_),
    .A2(_02363_),
    .B1(_02667_),
    .C1(_02668_),
    .Y(_02670_));
 sky130_fd_sc_hd__o211ai_2 _26777_ (.A1(net207),
    .A2(net204),
    .B1(_02669_),
    .C1(_02670_),
    .Y(_02671_));
 sky130_fd_sc_hd__o211ai_1 _26778_ (.A1(net200),
    .A2(_02362_),
    .B1(_02379_),
    .C1(_02667_),
    .Y(_02672_));
 sky130_fd_sc_hd__o2111ai_1 _26779_ (.A1(_08314_),
    .A2(_02363_),
    .B1(_02664_),
    .C1(_02666_),
    .D1(_02668_),
    .Y(_02673_));
 sky130_fd_sc_hd__nand3_2 _26780_ (.A(_07233_),
    .B(_02672_),
    .C(_02673_),
    .Y(_02675_));
 sky130_fd_sc_hd__o21ai_4 _26781_ (.A1(_07233_),
    .A2(_02661_),
    .B1(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__inv_2 _26782_ (.A(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__o211a_1 _26783_ (.A1(_02662_),
    .A2(_07233_),
    .B1(_08314_),
    .C1(_02671_),
    .X(_02678_));
 sky130_fd_sc_hd__o211ai_4 _26784_ (.A1(_02662_),
    .A2(_07233_),
    .B1(_08314_),
    .C1(_02671_),
    .Y(_02679_));
 sky130_fd_sc_hd__o211ai_4 _26785_ (.A1(_07233_),
    .A2(_02661_),
    .B1(net200),
    .C1(_02675_),
    .Y(_02680_));
 sky130_fd_sc_hd__nand2_1 _26786_ (.A(_02679_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__o2111a_1 _26787_ (.A1(_01438_),
    .A2(_01431_),
    .B1(_01437_),
    .C1(_01768_),
    .D1(_01770_),
    .X(_02682_));
 sky130_fd_sc_hd__o211a_1 _26788_ (.A1(_02058_),
    .A2(_02078_),
    .B1(_02682_),
    .C1(_02083_),
    .X(_02683_));
 sky130_fd_sc_hd__nand2_1 _26789_ (.A(_02386_),
    .B(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__o211ai_4 _26790_ (.A1(_02391_),
    .A2(_02385_),
    .B1(_02388_),
    .C1(_02684_),
    .Y(_02686_));
 sky130_fd_sc_hd__nand4_4 _26791_ (.A(_02683_),
    .B(_02388_),
    .C(_02386_),
    .D(_01445_),
    .Y(_02687_));
 sky130_fd_sc_hd__nand2_1 _26792_ (.A(_02686_),
    .B(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__a21oi_2 _26793_ (.A1(_02686_),
    .A2(_02687_),
    .B1(_02681_),
    .Y(_02689_));
 sky130_fd_sc_hd__a31o_1 _26794_ (.A1(_02681_),
    .A2(_02686_),
    .A3(_02687_),
    .B1(_07550_),
    .X(_02690_));
 sky130_fd_sc_hd__nand2_2 _26795_ (.A(_02676_),
    .B(_07550_),
    .Y(_02691_));
 sky130_fd_sc_hd__inv_2 _26796_ (.A(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__o211ai_4 _26797_ (.A1(_02676_),
    .A2(net197),
    .B1(_02687_),
    .C1(_02686_),
    .Y(_02693_));
 sky130_fd_sc_hd__nand4_4 _26798_ (.A(_02679_),
    .B(_02680_),
    .C(_02686_),
    .D(_02687_),
    .Y(_02694_));
 sky130_fd_sc_hd__a22o_1 _26799_ (.A1(_02679_),
    .A2(_02680_),
    .B1(_02686_),
    .B2(_02687_),
    .X(_02695_));
 sky130_fd_sc_hd__nand3_2 _26800_ (.A(_02695_),
    .B(_07548_),
    .C(_02694_),
    .Y(_02697_));
 sky130_fd_sc_hd__o221a_2 _26801_ (.A1(_07548_),
    .A2(_02676_),
    .B1(_02689_),
    .B2(_02690_),
    .C1(_07917_),
    .X(_02698_));
 sky130_fd_sc_hd__a211o_1 _26802_ (.A1(_02691_),
    .A2(_02697_),
    .B1(net183),
    .C1(net182),
    .X(_02699_));
 sky130_fd_sc_hd__a311oi_2 _26803_ (.A1(_02695_),
    .A2(_07548_),
    .A3(_02694_),
    .B1(_07936_),
    .C1(_02692_),
    .Y(_02700_));
 sky130_fd_sc_hd__nand3_4 _26804_ (.A(_02697_),
    .B(_07935_),
    .C(_02691_),
    .Y(_02701_));
 sky130_fd_sc_hd__o221ai_4 _26805_ (.A1(_07548_),
    .A2(_02676_),
    .B1(_02689_),
    .B2(_02690_),
    .C1(_07936_),
    .Y(_02702_));
 sky130_fd_sc_hd__a21oi_1 _26806_ (.A1(_02095_),
    .A2(_02398_),
    .B1(_02405_),
    .Y(_02703_));
 sky130_fd_sc_hd__o211a_1 _26807_ (.A1(net223),
    .A2(_02090_),
    .B1(_02398_),
    .C1(_02404_),
    .X(_02704_));
 sky130_fd_sc_hd__o22ai_2 _26808_ (.A1(_02383_),
    .A2(_02402_),
    .B1(_02405_),
    .B2(_02399_),
    .Y(_02705_));
 sky130_fd_sc_hd__a21boi_1 _26809_ (.A1(_02701_),
    .A2(_02702_),
    .B1_N(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__o2bb2ai_4 _26810_ (.A1_N(_02701_),
    .A2_N(_02702_),
    .B1(_02703_),
    .B2(_02403_),
    .Y(_02708_));
 sky130_fd_sc_hd__o211a_1 _26811_ (.A1(_02405_),
    .A2(_02704_),
    .B1(_02702_),
    .C1(_02701_),
    .X(_02709_));
 sky130_fd_sc_hd__o211ai_4 _26812_ (.A1(_02405_),
    .A2(_02704_),
    .B1(_02702_),
    .C1(_02701_),
    .Y(_02710_));
 sky130_fd_sc_hd__nand3_2 _26813_ (.A(_02708_),
    .B(_02710_),
    .C(net162),
    .Y(_02711_));
 sky130_fd_sc_hd__a311o_1 _26814_ (.A1(_02695_),
    .A2(_07548_),
    .A3(_02694_),
    .B1(net162),
    .C1(_02692_),
    .X(_02712_));
 sky130_fd_sc_hd__o22ai_1 _26815_ (.A1(net183),
    .A2(net182),
    .B1(_02706_),
    .B2(_02709_),
    .Y(_02713_));
 sky130_fd_sc_hd__a31oi_2 _26816_ (.A1(_02708_),
    .A2(_02710_),
    .A3(net162),
    .B1(_02698_),
    .Y(_02714_));
 sky130_fd_sc_hd__a31o_1 _26817_ (.A1(_02708_),
    .A2(_02710_),
    .A3(net162),
    .B1(_02698_),
    .X(_02715_));
 sky130_fd_sc_hd__o221ai_4 _26818_ (.A1(_06922_),
    .A2(_02101_),
    .B1(_02417_),
    .B2(_07246_),
    .C1(_02121_),
    .Y(_02716_));
 sky130_fd_sc_hd__a31oi_1 _26819_ (.A1(_02106_),
    .A2(_02121_),
    .A3(_02418_),
    .B1(_02419_),
    .Y(_02717_));
 sky130_fd_sc_hd__a311oi_4 _26820_ (.A1(_02708_),
    .A2(_02710_),
    .A3(net162),
    .B1(_02698_),
    .C1(_07565_),
    .Y(_02719_));
 sky130_fd_sc_hd__o211ai_4 _26821_ (.A1(_07560_),
    .A2(net217),
    .B1(_02699_),
    .C1(_02711_),
    .Y(_02720_));
 sky130_fd_sc_hd__a2bb2oi_2 _26822_ (.A1_N(net221),
    .A2_N(net219),
    .B1(_02699_),
    .B2(_02711_),
    .Y(_02721_));
 sky130_fd_sc_hd__o211ai_1 _26823_ (.A1(net221),
    .A2(net219),
    .B1(_02712_),
    .C1(_02713_),
    .Y(_02722_));
 sky130_fd_sc_hd__nor2_1 _26824_ (.A(_02719_),
    .B(_02721_),
    .Y(_02723_));
 sky130_fd_sc_hd__o2111ai_1 _26825_ (.A1(_02419_),
    .A2(_02424_),
    .B1(_02720_),
    .C1(_02722_),
    .D1(_02418_),
    .Y(_02724_));
 sky130_fd_sc_hd__o21ai_1 _26826_ (.A1(_02719_),
    .A2(_02721_),
    .B1(_02717_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand3_1 _26827_ (.A(_02724_),
    .B(_02725_),
    .C(net159),
    .Y(_02726_));
 sky130_fd_sc_hd__or3_1 _26828_ (.A(net181),
    .B(net179),
    .C(_02714_),
    .X(_02727_));
 sky130_fd_sc_hd__o211ai_2 _26829_ (.A1(_07564_),
    .A2(_02714_),
    .B1(_02716_),
    .C1(_02420_),
    .Y(_02728_));
 sky130_fd_sc_hd__o2bb2ai_1 _26830_ (.A1_N(_02420_),
    .A2_N(_02716_),
    .B1(_02719_),
    .B2(_02721_),
    .Y(_02730_));
 sky130_fd_sc_hd__o221ai_4 _26831_ (.A1(net181),
    .A2(net179),
    .B1(_02719_),
    .B2(_02728_),
    .C1(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__o21ai_2 _26832_ (.A1(net159),
    .A2(_02714_),
    .B1(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__inv_2 _26833_ (.A(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__o211a_1 _26834_ (.A1(_02715_),
    .A2(net159),
    .B1(net223),
    .C1(_02726_),
    .X(_02734_));
 sky130_fd_sc_hd__o211ai_4 _26835_ (.A1(_02715_),
    .A2(net159),
    .B1(net223),
    .C1(_02726_),
    .Y(_02735_));
 sky130_fd_sc_hd__nand3_4 _26836_ (.A(_02731_),
    .B(_07246_),
    .C(_02727_),
    .Y(_02736_));
 sky130_fd_sc_hd__nand2_2 _26837_ (.A(_02735_),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__o211ai_4 _26838_ (.A1(_02439_),
    .A2(_02431_),
    .B1(_02450_),
    .C1(_02447_),
    .Y(_02738_));
 sky130_fd_sc_hd__a31oi_2 _26839_ (.A1(_02441_),
    .A2(_02447_),
    .A3(_02450_),
    .B1(_02436_),
    .Y(_02739_));
 sky130_fd_sc_hd__o311a_2 _26840_ (.A1(_06918_),
    .A2(net249),
    .A3(_02432_),
    .B1(_02737_),
    .C1(_02738_),
    .X(_02741_));
 sky130_fd_sc_hd__o211ai_2 _26841_ (.A1(_06922_),
    .A2(_02432_),
    .B1(_02737_),
    .C1(_02738_),
    .Y(_02742_));
 sky130_fd_sc_hd__a21o_1 _26842_ (.A1(_02437_),
    .A2(_02738_),
    .B1(_02737_),
    .X(_02743_));
 sky130_fd_sc_hd__o22ai_4 _26843_ (.A1(net157),
    .A2(_08712_),
    .B1(_02737_),
    .B2(_02739_),
    .Y(_02744_));
 sky130_fd_sc_hd__nand3_2 _26844_ (.A(_02743_),
    .B(net149),
    .C(_02742_),
    .Y(_02745_));
 sky130_fd_sc_hd__and3_2 _26845_ (.A(_02732_),
    .B(_08713_),
    .C(_08710_),
    .X(_02746_));
 sky130_fd_sc_hd__inv_2 _26846_ (.A(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__o32a_2 _26847_ (.A1(net157),
    .A2(_08712_),
    .A3(_02733_),
    .B1(_02741_),
    .B2(_02744_),
    .X(_02748_));
 sky130_fd_sc_hd__o22ai_2 _26848_ (.A1(net149),
    .A2(_02733_),
    .B1(_02741_),
    .B2(_02744_),
    .Y(_02749_));
 sky130_fd_sc_hd__a311o_1 _26849_ (.A1(_02743_),
    .A2(net149),
    .A3(_02742_),
    .B1(_02746_),
    .C1(net146),
    .X(_02750_));
 sky130_fd_sc_hd__a22oi_4 _26850_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_02745_),
    .B2(_02747_),
    .Y(_02752_));
 sky130_fd_sc_hd__o21ai_4 _26851_ (.A1(_06914_),
    .A2(net250),
    .B1(_02749_),
    .Y(_02753_));
 sky130_fd_sc_hd__a31o_2 _26852_ (.A1(_02743_),
    .A2(net149),
    .A3(_02742_),
    .B1(net226),
    .X(_02754_));
 sky130_fd_sc_hd__o221a_1 _26853_ (.A1(net149),
    .A2(_02733_),
    .B1(_02741_),
    .B2(_02744_),
    .C1(_06922_),
    .X(_02755_));
 sky130_fd_sc_hd__o221ai_4 _26854_ (.A1(net149),
    .A2(_02733_),
    .B1(_02741_),
    .B2(_02744_),
    .C1(_06922_),
    .Y(_02756_));
 sky130_fd_sc_hd__a21oi_1 _26855_ (.A1(net233),
    .A2(_02460_),
    .B1(_02469_),
    .Y(_02757_));
 sky130_fd_sc_hd__nand2_1 _26856_ (.A(_02467_),
    .B(_02470_),
    .Y(_02758_));
 sky130_fd_sc_hd__a22oi_4 _26857_ (.A1(_02435_),
    .A2(_02463_),
    .B1(_02467_),
    .B2(_02470_),
    .Y(_02759_));
 sky130_fd_sc_hd__a22o_1 _26858_ (.A1(_02435_),
    .A2(_02463_),
    .B1(_02467_),
    .B2(_02470_),
    .X(_02760_));
 sky130_fd_sc_hd__o211ai_1 _26859_ (.A1(_02754_),
    .A2(_02746_),
    .B1(_02753_),
    .C1(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__o21ai_1 _26860_ (.A1(_02752_),
    .A2(_02755_),
    .B1(_02759_),
    .Y(_02763_));
 sky130_fd_sc_hd__o211ai_2 _26861_ (.A1(net148),
    .A2(net147),
    .B1(_02761_),
    .C1(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__a21oi_2 _26862_ (.A1(_02745_),
    .A2(_02747_),
    .B1(net146),
    .Y(_02765_));
 sky130_fd_sc_hd__o2bb2ai_4 _26863_ (.A1_N(_02753_),
    .A2_N(_02756_),
    .B1(_02757_),
    .B2(_02465_),
    .Y(_02766_));
 sky130_fd_sc_hd__o211ai_4 _26864_ (.A1(net233),
    .A2(_02460_),
    .B1(_02756_),
    .C1(_02758_),
    .Y(_02767_));
 sky130_fd_sc_hd__o211ai_2 _26865_ (.A1(_02746_),
    .A2(_02754_),
    .B1(_02753_),
    .C1(_02759_),
    .Y(_02768_));
 sky130_fd_sc_hd__o221ai_4 _26866_ (.A1(net148),
    .A2(net147),
    .B1(_02752_),
    .B2(_02767_),
    .C1(_02766_),
    .Y(_02769_));
 sky130_fd_sc_hd__a31o_1 _26867_ (.A1(net146),
    .A2(_02766_),
    .A3(_02768_),
    .B1(_02765_),
    .X(_02770_));
 sky130_fd_sc_hd__and3_1 _26868_ (.A(_02764_),
    .B(_09562_),
    .C(_02750_),
    .X(_02771_));
 sky130_fd_sc_hd__o21ai_2 _26869_ (.A1(_09559_),
    .A2(_09560_),
    .B1(_02770_),
    .Y(_02772_));
 sky130_fd_sc_hd__a311oi_4 _26870_ (.A1(net146),
    .A2(_02766_),
    .A3(_02768_),
    .B1(_02765_),
    .C1(net233),
    .Y(_02774_));
 sky130_fd_sc_hd__o211ai_4 _26871_ (.A1(net146),
    .A2(_02748_),
    .B1(net235),
    .C1(_02769_),
    .Y(_02775_));
 sky130_fd_sc_hd__o211ai_4 _26872_ (.A1(_06622_),
    .A2(_06624_),
    .B1(_02750_),
    .C1(_02764_),
    .Y(_02776_));
 sky130_fd_sc_hd__a21oi_1 _26873_ (.A1(_06315_),
    .A2(_02478_),
    .B1(_02481_),
    .Y(_02777_));
 sky130_fd_sc_hd__a31o_1 _26874_ (.A1(_06311_),
    .A2(_06313_),
    .A3(_02478_),
    .B1(_02481_),
    .X(_02778_));
 sky130_fd_sc_hd__o21ai_1 _26875_ (.A1(_02482_),
    .A2(_02483_),
    .B1(_02486_),
    .Y(_02779_));
 sky130_fd_sc_hd__a21oi_1 _26876_ (.A1(_02481_),
    .A2(_02484_),
    .B1(_02485_),
    .Y(_02780_));
 sky130_fd_sc_hd__a21oi_1 _26877_ (.A1(_02775_),
    .A2(_02776_),
    .B1(_02779_),
    .Y(_02781_));
 sky130_fd_sc_hd__o2bb2ai_2 _26878_ (.A1_N(_02775_),
    .A2_N(_02776_),
    .B1(_02777_),
    .B2(_02483_),
    .Y(_02782_));
 sky130_fd_sc_hd__o2111a_1 _26879_ (.A1(_06315_),
    .A2(_02478_),
    .B1(_02775_),
    .C1(_02776_),
    .D1(_02778_),
    .X(_02783_));
 sky130_fd_sc_hd__nand3_2 _26880_ (.A(_02779_),
    .B(_02776_),
    .C(_02775_),
    .Y(_02785_));
 sky130_fd_sc_hd__o211ai_2 _26881_ (.A1(net156),
    .A2(_09556_),
    .B1(_02782_),
    .C1(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__o22ai_2 _26882_ (.A1(net156),
    .A2(_09556_),
    .B1(_02781_),
    .B2(_02783_),
    .Y(_02787_));
 sky130_fd_sc_hd__o31a_2 _26883_ (.A1(_09562_),
    .A2(_02781_),
    .A3(_02783_),
    .B1(_02772_),
    .X(_02788_));
 sky130_fd_sc_hd__a31o_1 _26884_ (.A1(_09563_),
    .A2(_02782_),
    .A3(_02785_),
    .B1(_02771_),
    .X(_02789_));
 sky130_fd_sc_hd__o211ai_2 _26885_ (.A1(_05767_),
    .A2(_02180_),
    .B1(_02208_),
    .C1(_02498_),
    .Y(_02790_));
 sky130_fd_sc_hd__o2bb2ai_1 _26886_ (.A1_N(_02183_),
    .A2_N(_02208_),
    .B1(_06014_),
    .B2(_02495_),
    .Y(_02791_));
 sky130_fd_sc_hd__a31o_1 _26887_ (.A1(_09563_),
    .A2(_02782_),
    .A3(_02785_),
    .B1(_06315_),
    .X(_02792_));
 sky130_fd_sc_hd__a311oi_1 _26888_ (.A1(_09563_),
    .A2(_02782_),
    .A3(_02785_),
    .B1(_02771_),
    .C1(_06315_),
    .Y(_02793_));
 sky130_fd_sc_hd__o211ai_4 _26889_ (.A1(_06309_),
    .A2(_06312_),
    .B1(_02772_),
    .C1(_02786_),
    .Y(_02794_));
 sky130_fd_sc_hd__a2bb2oi_1 _26890_ (.A1_N(net284),
    .A2_N(net281),
    .B1(_02772_),
    .B2(_02786_),
    .Y(_02796_));
 sky130_fd_sc_hd__o221ai_4 _26891_ (.A1(net284),
    .A2(net281),
    .B1(_09563_),
    .B2(_02770_),
    .C1(_02787_),
    .Y(_02797_));
 sky130_fd_sc_hd__o2111ai_1 _26892_ (.A1(_02496_),
    .A2(_06013_),
    .B1(_02794_),
    .C1(_02791_),
    .D1(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__o2bb2ai_1 _26893_ (.A1_N(_02498_),
    .A2_N(_02791_),
    .B1(_02793_),
    .B2(_02796_),
    .Y(_02799_));
 sky130_fd_sc_hd__o211ai_2 _26894_ (.A1(net142),
    .A2(_09573_),
    .B1(_02798_),
    .C1(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__o2111ai_1 _26895_ (.A1(_06014_),
    .A2(_02495_),
    .B1(_02790_),
    .C1(_02794_),
    .D1(_02797_),
    .Y(_02801_));
 sky130_fd_sc_hd__o2bb2ai_1 _26896_ (.A1_N(_02501_),
    .A2_N(_02790_),
    .B1(_02793_),
    .B2(_02796_),
    .Y(_02802_));
 sky130_fd_sc_hd__o211ai_2 _26897_ (.A1(net142),
    .A2(_09573_),
    .B1(_02801_),
    .C1(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__o31a_2 _26898_ (.A1(net142),
    .A2(_09573_),
    .A3(_02788_),
    .B1(_02803_),
    .X(_02804_));
 sky130_fd_sc_hd__o21ai_1 _26899_ (.A1(_10477_),
    .A2(_10478_),
    .B1(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__o211ai_4 _26900_ (.A1(net132),
    .A2(_02789_),
    .B1(_02800_),
    .C1(_06014_),
    .Y(_02807_));
 sky130_fd_sc_hd__o221a_1 _26901_ (.A1(net285),
    .A2(_06012_),
    .B1(net132),
    .B2(_02788_),
    .C1(_02803_),
    .X(_02808_));
 sky130_fd_sc_hd__o221ai_2 _26902_ (.A1(net285),
    .A2(_06012_),
    .B1(net132),
    .B2(_02788_),
    .C1(_02803_),
    .Y(_02809_));
 sky130_fd_sc_hd__nand2_1 _26903_ (.A(_02807_),
    .B(_02809_),
    .Y(_02810_));
 sky130_fd_sc_hd__a31o_1 _26904_ (.A1(_02514_),
    .A2(_02519_),
    .A3(_02522_),
    .B1(_02511_),
    .X(_02811_));
 sky130_fd_sc_hd__a31oi_4 _26905_ (.A1(_02514_),
    .A2(_02519_),
    .A3(_02522_),
    .B1(_02511_),
    .Y(_02812_));
 sky130_fd_sc_hd__and4_1 _26906_ (.A(_02512_),
    .B(_02525_),
    .C(_02807_),
    .D(_02809_),
    .X(_02813_));
 sky130_fd_sc_hd__o2bb2ai_1 _26907_ (.A1_N(_02810_),
    .A2_N(_02811_),
    .B1(net141),
    .B2(net140),
    .Y(_02814_));
 sky130_fd_sc_hd__nand2_1 _26908_ (.A(_02810_),
    .B(_02812_),
    .Y(_02815_));
 sky130_fd_sc_hd__a21o_1 _26909_ (.A1(_02512_),
    .A2(_02525_),
    .B1(_02810_),
    .X(_02816_));
 sky130_fd_sc_hd__o211ai_4 _26910_ (.A1(net141),
    .A2(net140),
    .B1(_02815_),
    .C1(_02816_),
    .Y(_02818_));
 sky130_fd_sc_hd__o21ai_4 _26911_ (.A1(net131),
    .A2(_02804_),
    .B1(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__o211ai_4 _26912_ (.A1(_02813_),
    .A2(_02814_),
    .B1(_05768_),
    .C1(_02805_),
    .Y(_02820_));
 sky130_fd_sc_hd__inv_2 _26913_ (.A(_02820_),
    .Y(_02821_));
 sky130_fd_sc_hd__o221ai_4 _26914_ (.A1(_05765_),
    .A2(net288),
    .B1(net131),
    .B2(_02804_),
    .C1(_02818_),
    .Y(_02822_));
 sky130_fd_sc_hd__nand2_1 _26915_ (.A(_02820_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__a21oi_1 _26916_ (.A1(_01900_),
    .A2(_04238_),
    .B1(_01569_),
    .Y(_02824_));
 sky130_fd_sc_hd__o2111a_1 _26917_ (.A1(_04238_),
    .A2(_01900_),
    .B1(_02824_),
    .C1(_02229_),
    .D1(_02227_),
    .X(_02825_));
 sky130_fd_sc_hd__nand2_1 _26918_ (.A(_02535_),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__o211ai_4 _26919_ (.A1(_02533_),
    .A2(_02534_),
    .B1(_02537_),
    .C1(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__nand4_4 _26920_ (.A(_02825_),
    .B(_02537_),
    .C(_02535_),
    .D(_01575_),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _26921_ (.A(_02827_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__nand3_1 _26922_ (.A(_02823_),
    .B(_02827_),
    .C(_02829_),
    .Y(_02831_));
 sky130_fd_sc_hd__a21o_1 _26923_ (.A1(_02827_),
    .A2(_02829_),
    .B1(_02823_),
    .X(_02832_));
 sky130_fd_sc_hd__o211ai_2 _26924_ (.A1(net137),
    .A2(net135),
    .B1(_02831_),
    .C1(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__or3b_2 _26925_ (.A(net137),
    .B(net135),
    .C_N(_02819_),
    .X(_02834_));
 sky130_fd_sc_hd__a22oi_1 _26926_ (.A1(_02820_),
    .A2(_02822_),
    .B1(_02827_),
    .B2(_02829_),
    .Y(_02835_));
 sky130_fd_sc_hd__a22o_1 _26927_ (.A1(_02820_),
    .A2(_02822_),
    .B1(_02827_),
    .B2(_02829_),
    .X(_02836_));
 sky130_fd_sc_hd__o211ai_4 _26928_ (.A1(_02819_),
    .A2(_05768_),
    .B1(_02829_),
    .C1(_02827_),
    .Y(_02837_));
 sky130_fd_sc_hd__o2111a_1 _26929_ (.A1(_05768_),
    .A2(_02819_),
    .B1(_02820_),
    .C1(_02827_),
    .D1(_02829_),
    .X(_02838_));
 sky130_fd_sc_hd__o221ai_4 _26930_ (.A1(net137),
    .A2(net135),
    .B1(_02821_),
    .B2(_02837_),
    .C1(_02836_),
    .Y(_02840_));
 sky130_fd_sc_hd__o21a_1 _26931_ (.A1(_10954_),
    .A2(_02819_),
    .B1(_02833_),
    .X(_02841_));
 sky130_fd_sc_hd__o311a_1 _26932_ (.A1(_10953_),
    .A2(_02835_),
    .A3(_02838_),
    .B1(_02834_),
    .C1(_05507_),
    .X(_02842_));
 sky130_fd_sc_hd__o211ai_4 _26933_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_02834_),
    .C1(_02840_),
    .Y(_02843_));
 sky130_fd_sc_hd__o211ai_4 _26934_ (.A1(_02819_),
    .A2(_10954_),
    .B1(_05508_),
    .C1(_02833_),
    .Y(_02844_));
 sky130_fd_sc_hd__a21o_1 _26935_ (.A1(_02549_),
    .A2(_02547_),
    .B1(_02544_),
    .X(_02845_));
 sky130_fd_sc_hd__a21oi_1 _26936_ (.A1(_02549_),
    .A2(_02547_),
    .B1(_02544_),
    .Y(_02846_));
 sky130_fd_sc_hd__a21o_1 _26937_ (.A1(_02843_),
    .A2(_02844_),
    .B1(_02845_),
    .X(_02847_));
 sky130_fd_sc_hd__a31oi_2 _26938_ (.A1(_02845_),
    .A2(_02844_),
    .A3(_02843_),
    .B1(_11464_),
    .Y(_02848_));
 sky130_fd_sc_hd__a22oi_2 _26939_ (.A1(_11464_),
    .A2(_02841_),
    .B1(_02847_),
    .B2(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__a21oi_2 _26940_ (.A1(_05243_),
    .A2(_05245_),
    .B1(_02849_),
    .Y(_02851_));
 sky130_fd_sc_hd__a221oi_2 _26941_ (.A1(_11464_),
    .A2(_02841_),
    .B1(_02847_),
    .B2(_02848_),
    .C1(_05249_),
    .Y(_02852_));
 sky130_fd_sc_hd__a221o_1 _26942_ (.A1(_11464_),
    .A2(_02841_),
    .B1(_02847_),
    .B2(_02848_),
    .C1(_05249_),
    .X(_02853_));
 sky130_fd_sc_hd__o21ai_1 _26943_ (.A1(_02553_),
    .A2(_02557_),
    .B1(_02556_),
    .Y(_02854_));
 sky130_fd_sc_hd__o221ai_1 _26944_ (.A1(_02557_),
    .A2(_02553_),
    .B1(_02852_),
    .B2(_02851_),
    .C1(_02556_),
    .Y(_02855_));
 sky130_fd_sc_hd__a21bo_1 _26945_ (.A1(_02855_),
    .A2(net133),
    .B1_N(_02849_),
    .X(_02856_));
 sky130_fd_sc_hd__a21oi_1 _26946_ (.A1(_05119_),
    .A2(_02562_),
    .B1(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__and3_1 _26947_ (.A(_05119_),
    .B(_02562_),
    .C(_02856_),
    .X(_02858_));
 sky130_fd_sc_hd__nor2_1 _26948_ (.A(_02857_),
    .B(_02858_),
    .Y(net104));
 sky130_fd_sc_hd__or3_1 _26949_ (.A(_02260_),
    .B(_02559_),
    .C(_02856_),
    .X(_02859_));
 sky130_fd_sc_hd__and4_1 _26950_ (.A(_01784_),
    .B(_01786_),
    .C(_02092_),
    .D(_02095_),
    .X(_02861_));
 sky130_fd_sc_hd__o211a_1 _26951_ (.A1(_02383_),
    .A2(_02402_),
    .B1(_02861_),
    .C1(_02406_),
    .X(_02862_));
 sky130_fd_sc_hd__nand3_1 _26952_ (.A(_02701_),
    .B(_02861_),
    .C(_02407_),
    .Y(_02863_));
 sky130_fd_sc_hd__o211ai_4 _26953_ (.A1(_02705_),
    .A2(_02700_),
    .B1(_02702_),
    .C1(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__nand4_4 _26954_ (.A(_02862_),
    .B(_02702_),
    .C(_02701_),
    .D(_01795_),
    .Y(_02865_));
 sky130_fd_sc_hd__and2_1 _26955_ (.A(_02864_),
    .B(_02865_),
    .X(_02866_));
 sky130_fd_sc_hd__a31o_2 _26956_ (.A1(_11471_),
    .A2(_02568_),
    .A3(_02573_),
    .B1(_05754_),
    .X(_02867_));
 sky130_fd_sc_hd__a311o_1 _26957_ (.A1(_11471_),
    .A2(_02568_),
    .A3(_02573_),
    .B1(net240),
    .C1(_05754_),
    .X(_02868_));
 sky130_fd_sc_hd__o311a_1 _26958_ (.A1(_11470_),
    .A2(_02567_),
    .A3(_02572_),
    .B1(_10971_),
    .C1(_05752_),
    .X(_02869_));
 sky130_fd_sc_hd__o21a_1 _26959_ (.A1(_10965_),
    .A2(_10967_),
    .B1(_02867_),
    .X(_02870_));
 sky130_fd_sc_hd__nor2_1 _26960_ (.A(_02869_),
    .B(_02870_),
    .Y(_02872_));
 sky130_fd_sc_hd__o221ai_2 _26961_ (.A1(_02293_),
    .A2(net153),
    .B1(net150),
    .B2(_02580_),
    .C1(_02591_),
    .Y(_02873_));
 sky130_fd_sc_hd__a22oi_2 _26962_ (.A1(net150),
    .A2(_02580_),
    .B1(_02591_),
    .B2(_02294_),
    .Y(_02874_));
 sky130_fd_sc_hd__nand3_2 _26963_ (.A(_02585_),
    .B(_02873_),
    .C(_02872_),
    .Y(_02875_));
 sky130_fd_sc_hd__o311ai_4 _26964_ (.A1(_02582_),
    .A2(_02872_),
    .A3(_02874_),
    .B1(_02875_),
    .C1(net240),
    .Y(_02876_));
 sky130_fd_sc_hd__o31a_1 _26965_ (.A1(net260),
    .A2(net255),
    .A3(_02867_),
    .B1(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__o21ai_4 _26966_ (.A1(net240),
    .A2(_02867_),
    .B1(_02876_),
    .Y(_02878_));
 sky130_fd_sc_hd__a2bb2oi_2 _26967_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_02868_),
    .B2(_02876_),
    .Y(_02879_));
 sky130_fd_sc_hd__a2bb2o_2 _26968_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_02868_),
    .B2(_02876_),
    .X(_02880_));
 sky130_fd_sc_hd__o211a_2 _26969_ (.A1(net240),
    .A2(_02867_),
    .B1(net150),
    .C1(_02876_),
    .X(_02881_));
 sky130_fd_sc_hd__o211ai_1 _26970_ (.A1(net240),
    .A2(_02867_),
    .B1(net150),
    .C1(_02876_),
    .Y(_02883_));
 sky130_fd_sc_hd__nor2_1 _26971_ (.A(_02879_),
    .B(_02881_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_1 _26972_ (.A(_02880_),
    .B(_02883_),
    .Y(_02885_));
 sky130_fd_sc_hd__o21a_1 _26973_ (.A1(net151),
    .A2(_02600_),
    .B1(_02614_),
    .X(_02886_));
 sky130_fd_sc_hd__o21ai_1 _26974_ (.A1(net151),
    .A2(_02600_),
    .B1(_02614_),
    .Y(_02887_));
 sky130_fd_sc_hd__a22oi_4 _26975_ (.A1(net151),
    .A2(_02600_),
    .B1(_02886_),
    .B2(_02613_),
    .Y(_02888_));
 sky130_fd_sc_hd__o211a_1 _26976_ (.A1(net153),
    .A2(_02601_),
    .B1(_02617_),
    .C1(_02884_),
    .X(_02889_));
 sky130_fd_sc_hd__o21ai_2 _26977_ (.A1(_02884_),
    .A2(_02888_),
    .B1(_06293_),
    .Y(_02890_));
 sky130_fd_sc_hd__or3_1 _26978_ (.A(net239),
    .B(_06292_),
    .C(_02877_),
    .X(_02891_));
 sky130_fd_sc_hd__o221ai_4 _26979_ (.A1(net153),
    .A2(_02601_),
    .B1(_02879_),
    .B2(_02881_),
    .C1(_02617_),
    .Y(_02892_));
 sky130_fd_sc_hd__o211ai_4 _26980_ (.A1(_02885_),
    .A2(_02888_),
    .B1(_02892_),
    .C1(_06293_),
    .Y(_02894_));
 sky130_fd_sc_hd__o21ai_4 _26981_ (.A1(_06293_),
    .A2(_02877_),
    .B1(_02894_),
    .Y(_02895_));
 sky130_fd_sc_hd__inv_2 _26982_ (.A(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__o221ai_4 _26983_ (.A1(_06293_),
    .A2(_02878_),
    .B1(_02889_),
    .B2(_02890_),
    .C1(net151),
    .Y(_02897_));
 sky130_fd_sc_hd__o211ai_2 _26984_ (.A1(net167),
    .A2(_10024_),
    .B1(_02891_),
    .C1(_02894_),
    .Y(_02898_));
 sky130_fd_sc_hd__nand2_1 _26985_ (.A(_02897_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__and3_1 _26986_ (.A(_02017_),
    .B(_02019_),
    .C(_01714_),
    .X(_02900_));
 sky130_fd_sc_hd__o211ai_1 _26987_ (.A1(_02318_),
    .A2(_02339_),
    .B1(_02900_),
    .C1(_02343_),
    .Y(_02901_));
 sky130_fd_sc_hd__a31oi_1 _26988_ (.A1(_02620_),
    .A2(net172),
    .A3(_02602_),
    .B1(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__a31o_1 _26989_ (.A1(_02620_),
    .A2(net172),
    .A3(_02602_),
    .B1(_02901_),
    .X(_02903_));
 sky130_fd_sc_hd__a211oi_1 _26990_ (.A1(_02634_),
    .A2(_02628_),
    .B1(_02629_),
    .C1(_02902_),
    .Y(_02905_));
 sky130_fd_sc_hd__o211ai_4 _26991_ (.A1(_02635_),
    .A2(_02627_),
    .B1(_02631_),
    .C1(_02903_),
    .Y(_02906_));
 sky130_fd_sc_hd__nand4_1 _26992_ (.A(_02900_),
    .B(_02343_),
    .C(_02341_),
    .D(_01728_),
    .Y(_02907_));
 sky130_fd_sc_hd__nand3b_4 _26993_ (.A_N(_02907_),
    .B(_02631_),
    .C(_02628_),
    .Y(_02908_));
 sky130_fd_sc_hd__nand3_1 _26994_ (.A(_02899_),
    .B(_02906_),
    .C(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__a21o_1 _26995_ (.A1(_02906_),
    .A2(_02908_),
    .B1(_02899_),
    .X(_02910_));
 sky130_fd_sc_hd__nand4_2 _26996_ (.A(_02897_),
    .B(_02898_),
    .C(_02906_),
    .D(_02908_),
    .Y(_02911_));
 sky130_fd_sc_hd__a22o_1 _26997_ (.A1(_02897_),
    .A2(_02898_),
    .B1(_02906_),
    .B2(_02908_),
    .X(_02912_));
 sky130_fd_sc_hd__nand3_2 _26998_ (.A(_02912_),
    .B(net209),
    .C(_02911_),
    .Y(_02913_));
 sky130_fd_sc_hd__o221a_1 _26999_ (.A1(_06293_),
    .A2(_02878_),
    .B1(_02889_),
    .B2(_02890_),
    .C1(_06613_),
    .X(_02914_));
 sky130_fd_sc_hd__a211o_1 _27000_ (.A1(_02891_),
    .A2(_02894_),
    .B1(net238),
    .C1(net236),
    .X(_02916_));
 sky130_fd_sc_hd__or3_1 _27001_ (.A(net238),
    .B(net236),
    .C(_02895_),
    .X(_02917_));
 sky130_fd_sc_hd__o211ai_2 _27002_ (.A1(net238),
    .A2(net236),
    .B1(_02909_),
    .C1(_02910_),
    .Y(_02918_));
 sky130_fd_sc_hd__o221a_2 _27003_ (.A1(_06897_),
    .A2(_06898_),
    .B1(_02895_),
    .B2(net209),
    .C1(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__a211o_1 _27004_ (.A1(_02913_),
    .A2(_02916_),
    .B1(net229),
    .C1(net228),
    .X(_02920_));
 sky130_fd_sc_hd__a311oi_4 _27005_ (.A1(_02912_),
    .A2(net209),
    .A3(_02911_),
    .B1(_02914_),
    .C1(net171),
    .Y(_02921_));
 sky130_fd_sc_hd__nand3_4 _27006_ (.A(_02913_),
    .B(_02916_),
    .C(net172),
    .Y(_02922_));
 sky130_fd_sc_hd__o211ai_4 _27007_ (.A1(net189),
    .A2(net188),
    .B1(_02917_),
    .C1(_02918_),
    .Y(_02923_));
 sky130_fd_sc_hd__o211a_1 _27008_ (.A1(_02359_),
    .A2(_02353_),
    .B1(_02352_),
    .C1(_02653_),
    .X(_02924_));
 sky130_fd_sc_hd__o22ai_4 _27009_ (.A1(_02625_),
    .A2(_02648_),
    .B1(_02651_),
    .B2(_02646_),
    .Y(_02925_));
 sky130_fd_sc_hd__o2bb2ai_4 _27010_ (.A1_N(_02922_),
    .A2_N(_02923_),
    .B1(_02924_),
    .B2(_02649_),
    .Y(_02927_));
 sky130_fd_sc_hd__nand3b_4 _27011_ (.A_N(_02925_),
    .B(_02923_),
    .C(_02922_),
    .Y(_02928_));
 sky130_fd_sc_hd__nand3_1 _27012_ (.A(_02927_),
    .B(_02928_),
    .C(_06903_),
    .Y(_02929_));
 sky130_fd_sc_hd__a31oi_4 _27013_ (.A1(_02927_),
    .A2(_02928_),
    .A3(_06903_),
    .B1(_02919_),
    .Y(_02930_));
 sky130_fd_sc_hd__a311o_2 _27014_ (.A1(_02927_),
    .A2(_02928_),
    .A3(_06903_),
    .B1(_07233_),
    .C1(_02919_),
    .X(_02931_));
 sky130_fd_sc_hd__o221ai_1 _27015_ (.A1(net178),
    .A2(_02661_),
    .B1(_02362_),
    .B2(net200),
    .C1(_02379_),
    .Y(_02932_));
 sky130_fd_sc_hd__a31oi_2 _27016_ (.A1(_02368_),
    .A2(_02379_),
    .A3(_02664_),
    .B1(_02665_),
    .Y(_02933_));
 sky130_fd_sc_hd__o21ai_1 _27017_ (.A1(_08731_),
    .A2(_02662_),
    .B1(_02932_),
    .Y(_02934_));
 sky130_fd_sc_hd__a311oi_4 _27018_ (.A1(_02927_),
    .A2(_02928_),
    .A3(_06903_),
    .B1(_09140_),
    .C1(_02919_),
    .Y(_02935_));
 sky130_fd_sc_hd__nand3_1 _27019_ (.A(_02929_),
    .B(_09139_),
    .C(_02920_),
    .Y(_02936_));
 sky130_fd_sc_hd__a2bb2oi_2 _27020_ (.A1_N(net194),
    .A2_N(net191),
    .B1(_02920_),
    .B2(_02929_),
    .Y(_02938_));
 sky130_fd_sc_hd__a2bb2o_1 _27021_ (.A1_N(net194),
    .A2_N(net191),
    .B1(_02920_),
    .B2(_02929_),
    .X(_02939_));
 sky130_fd_sc_hd__nor2_1 _27022_ (.A(_02935_),
    .B(_02938_),
    .Y(_02940_));
 sky130_fd_sc_hd__nand3_1 _27023_ (.A(_02934_),
    .B(_02936_),
    .C(_02939_),
    .Y(_02941_));
 sky130_fd_sc_hd__o21ai_1 _27024_ (.A1(_02935_),
    .A2(_02938_),
    .B1(_02933_),
    .Y(_02942_));
 sky130_fd_sc_hd__o211ai_4 _27025_ (.A1(net207),
    .A2(net204),
    .B1(_02941_),
    .C1(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__o21ai_1 _27026_ (.A1(_09139_),
    .A2(_02930_),
    .B1(_02933_),
    .Y(_02944_));
 sky130_fd_sc_hd__o21ai_1 _27027_ (.A1(_02935_),
    .A2(_02938_),
    .B1(_02934_),
    .Y(_02945_));
 sky130_fd_sc_hd__o221ai_4 _27028_ (.A1(net207),
    .A2(net204),
    .B1(_02935_),
    .B2(_02944_),
    .C1(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__o21ai_2 _27029_ (.A1(_07233_),
    .A2(_02930_),
    .B1(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__nand2_2 _27030_ (.A(_02931_),
    .B(_02943_),
    .Y(_02949_));
 sky130_fd_sc_hd__o311a_1 _27031_ (.A1(net207),
    .A2(net204),
    .A3(_02930_),
    .B1(_02946_),
    .C1(_07550_),
    .X(_02950_));
 sky130_fd_sc_hd__o211a_1 _27032_ (.A1(_08724_),
    .A2(net196),
    .B1(_02931_),
    .C1(_02943_),
    .X(_02951_));
 sky130_fd_sc_hd__o211ai_4 _27033_ (.A1(_08724_),
    .A2(net196),
    .B1(_02931_),
    .C1(_02943_),
    .Y(_02952_));
 sky130_fd_sc_hd__o311a_1 _27034_ (.A1(net207),
    .A2(net204),
    .A3(_02930_),
    .B1(net178),
    .C1(_02946_),
    .X(_02953_));
 sky130_fd_sc_hd__o211ai_4 _27035_ (.A1(_07233_),
    .A2(_02930_),
    .B1(net178),
    .C1(_02946_),
    .Y(_02954_));
 sky130_fd_sc_hd__nand2_1 _27036_ (.A(_02952_),
    .B(_02954_),
    .Y(_02955_));
 sky130_fd_sc_hd__a31oi_1 _27037_ (.A1(_02680_),
    .A2(_02686_),
    .A3(_02687_),
    .B1(_02678_),
    .Y(_02956_));
 sky130_fd_sc_hd__o2bb2a_1 _27038_ (.A1_N(_02679_),
    .A2_N(_02693_),
    .B1(_02951_),
    .B2(_02953_),
    .X(_02957_));
 sky130_fd_sc_hd__a22o_1 _27039_ (.A1(_02679_),
    .A2(_02693_),
    .B1(_02952_),
    .B2(_02954_),
    .X(_02958_));
 sky130_fd_sc_hd__o2111ai_2 _27040_ (.A1(net201),
    .A2(_02677_),
    .B1(_02693_),
    .C1(_02952_),
    .D1(_02954_),
    .Y(_02960_));
 sky130_fd_sc_hd__a41o_1 _27041_ (.A1(_02679_),
    .A2(_02693_),
    .A3(_02952_),
    .A4(_02954_),
    .B1(_07550_),
    .X(_02961_));
 sky130_fd_sc_hd__o221a_1 _27042_ (.A1(_02677_),
    .A2(net200),
    .B1(_02953_),
    .B2(_02951_),
    .C1(_02694_),
    .X(_02962_));
 sky130_fd_sc_hd__o21ai_2 _27043_ (.A1(_02955_),
    .A2(_02956_),
    .B1(_07548_),
    .Y(_02963_));
 sky130_fd_sc_hd__o22a_1 _27044_ (.A1(_07548_),
    .A2(_02947_),
    .B1(_02961_),
    .B2(_02957_),
    .X(_02964_));
 sky130_fd_sc_hd__a31o_1 _27045_ (.A1(_02958_),
    .A2(_02960_),
    .A3(_07548_),
    .B1(_02950_),
    .X(_02965_));
 sky130_fd_sc_hd__o221a_1 _27046_ (.A1(_07548_),
    .A2(_02947_),
    .B1(_02961_),
    .B2(_02957_),
    .C1(net197),
    .X(_02966_));
 sky130_fd_sc_hd__a311o_2 _27047_ (.A1(_02958_),
    .A2(_02960_),
    .A3(_07548_),
    .B1(net201),
    .C1(_02950_),
    .X(_02967_));
 sky130_fd_sc_hd__o221a_1 _27048_ (.A1(_07548_),
    .A2(_02949_),
    .B1(_02963_),
    .B2(_02962_),
    .C1(net200),
    .X(_02968_));
 sky130_fd_sc_hd__o221ai_4 _27049_ (.A1(_07548_),
    .A2(_02949_),
    .B1(_02963_),
    .B2(_02962_),
    .C1(net201),
    .Y(_02969_));
 sky130_fd_sc_hd__o2bb2ai_4 _27050_ (.A1_N(_02864_),
    .A2_N(_02865_),
    .B1(_02966_),
    .B2(_02968_),
    .Y(_02971_));
 sky130_fd_sc_hd__nand4_4 _27051_ (.A(_02864_),
    .B(_02865_),
    .C(_02967_),
    .D(_02969_),
    .Y(_02972_));
 sky130_fd_sc_hd__nand3_2 _27052_ (.A(_02971_),
    .B(_02972_),
    .C(net162),
    .Y(_02973_));
 sky130_fd_sc_hd__o221a_2 _27053_ (.A1(_07548_),
    .A2(_02947_),
    .B1(_02961_),
    .B2(_02957_),
    .C1(_07917_),
    .X(_02974_));
 sky130_fd_sc_hd__a311o_2 _27054_ (.A1(_02958_),
    .A2(_02960_),
    .A3(_07548_),
    .B1(_07916_),
    .C1(_02950_),
    .X(_02975_));
 sky130_fd_sc_hd__a31oi_1 _27055_ (.A1(_02971_),
    .A2(_02972_),
    .A3(net162),
    .B1(_02974_),
    .Y(_02976_));
 sky130_fd_sc_hd__a21oi_2 _27056_ (.A1(_02973_),
    .A2(_02975_),
    .B1(net159),
    .Y(_02977_));
 sky130_fd_sc_hd__or3_2 _27057_ (.A(net181),
    .B(net179),
    .C(_02976_),
    .X(_02978_));
 sky130_fd_sc_hd__a31o_1 _27058_ (.A1(_02971_),
    .A2(_02972_),
    .A3(net162),
    .B1(_07936_),
    .X(_02979_));
 sky130_fd_sc_hd__a311oi_4 _27059_ (.A1(_02971_),
    .A2(_02972_),
    .A3(net162),
    .B1(_02974_),
    .C1(_07936_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand3_2 _27060_ (.A(_02973_),
    .B(_02975_),
    .C(_07935_),
    .Y(_02982_));
 sky130_fd_sc_hd__a22oi_2 _27061_ (.A1(_07929_),
    .A2(_07932_),
    .B1(_02973_),
    .B2(_02975_),
    .Y(_02983_));
 sky130_fd_sc_hd__a22o_2 _27062_ (.A1(_07929_),
    .A2(_07932_),
    .B1(_02973_),
    .B2(_02975_),
    .X(_02984_));
 sky130_fd_sc_hd__a31o_1 _27063_ (.A1(_02420_),
    .A2(_02716_),
    .A3(_02720_),
    .B1(_02721_),
    .X(_02985_));
 sky130_fd_sc_hd__a31oi_2 _27064_ (.A1(_02420_),
    .A2(_02716_),
    .A3(_02720_),
    .B1(_02721_),
    .Y(_02986_));
 sky130_fd_sc_hd__o21bai_4 _27065_ (.A1(_02980_),
    .A2(_02983_),
    .B1_N(_02985_),
    .Y(_02987_));
 sky130_fd_sc_hd__o21ai_1 _27066_ (.A1(_07935_),
    .A2(_02976_),
    .B1(_02985_),
    .Y(_02988_));
 sky130_fd_sc_hd__o211ai_2 _27067_ (.A1(_02974_),
    .A2(_02979_),
    .B1(_02985_),
    .C1(_02984_),
    .Y(_02989_));
 sky130_fd_sc_hd__o211ai_4 _27068_ (.A1(_02980_),
    .A2(_02988_),
    .B1(net159),
    .C1(_02987_),
    .Y(_02990_));
 sky130_fd_sc_hd__a31o_2 _27069_ (.A1(_02987_),
    .A2(_02989_),
    .A3(net159),
    .B1(_02977_),
    .X(_02991_));
 sky130_fd_sc_hd__o211ai_4 _27070_ (.A1(_06922_),
    .A2(_02432_),
    .B1(_02735_),
    .C1(_02738_),
    .Y(_02993_));
 sky130_fd_sc_hd__a2bb2oi_1 _27071_ (.A1_N(_02732_),
    .A2_N(net223),
    .B1(_02437_),
    .B2(_02738_),
    .Y(_02994_));
 sky130_fd_sc_hd__o21ai_1 _27072_ (.A1(net223),
    .A2(_02732_),
    .B1(_02993_),
    .Y(_02995_));
 sky130_fd_sc_hd__a311oi_4 _27073_ (.A1(_02987_),
    .A2(_02989_),
    .A3(net159),
    .B1(_02977_),
    .C1(_07565_),
    .Y(_02996_));
 sky130_fd_sc_hd__nand3_2 _27074_ (.A(_02990_),
    .B(_07564_),
    .C(_02978_),
    .Y(_02997_));
 sky130_fd_sc_hd__a22oi_4 _27075_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_02978_),
    .B2(_02990_),
    .Y(_02998_));
 sky130_fd_sc_hd__a22o_1 _27076_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_02978_),
    .B2(_02990_),
    .X(_02999_));
 sky130_fd_sc_hd__nand3_1 _27077_ (.A(_02995_),
    .B(_02997_),
    .C(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__o22ai_1 _27078_ (.A1(_02734_),
    .A2(_02994_),
    .B1(_02996_),
    .B2(_02998_),
    .Y(_03001_));
 sky130_fd_sc_hd__nand3_2 _27079_ (.A(_03000_),
    .B(_03001_),
    .C(net149),
    .Y(_03002_));
 sky130_fd_sc_hd__and3_1 _27080_ (.A(_08710_),
    .B(_08713_),
    .C(_02991_),
    .X(_03004_));
 sky130_fd_sc_hd__a22o_1 _27081_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_02978_),
    .B2(_02990_),
    .X(_03005_));
 sky130_fd_sc_hd__o211ai_2 _27082_ (.A1(_02734_),
    .A2(_02994_),
    .B1(_02997_),
    .C1(_02999_),
    .Y(_03006_));
 sky130_fd_sc_hd__o2bb2ai_1 _27083_ (.A1_N(_02736_),
    .A2_N(_02993_),
    .B1(_02996_),
    .B2(_02998_),
    .Y(_03007_));
 sky130_fd_sc_hd__o211ai_2 _27084_ (.A1(net157),
    .A2(_08712_),
    .B1(_03006_),
    .C1(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__a31o_1 _27085_ (.A1(_03006_),
    .A2(_03007_),
    .A3(net149),
    .B1(_03004_),
    .X(_03009_));
 sky130_fd_sc_hd__o21ai_4 _27086_ (.A1(net149),
    .A2(_02991_),
    .B1(_03002_),
    .Y(_03010_));
 sky130_fd_sc_hd__o211ai_4 _27087_ (.A1(_02991_),
    .A2(net149),
    .B1(net223),
    .C1(_03002_),
    .Y(_03011_));
 sky130_fd_sc_hd__a31o_1 _27088_ (.A1(_03006_),
    .A2(_03007_),
    .A3(net149),
    .B1(net223),
    .X(_03012_));
 sky130_fd_sc_hd__o211ai_4 _27089_ (.A1(_07244_),
    .A2(net247),
    .B1(_03005_),
    .C1(_03008_),
    .Y(_03013_));
 sky130_fd_sc_hd__a22oi_1 _27090_ (.A1(net226),
    .A2(_02749_),
    .B1(_02758_),
    .B2(_02464_),
    .Y(_03015_));
 sky130_fd_sc_hd__a31o_1 _27091_ (.A1(_02464_),
    .A2(_02756_),
    .A3(_02758_),
    .B1(_02752_),
    .X(_03016_));
 sky130_fd_sc_hd__o22ai_2 _27092_ (.A1(_02754_),
    .A2(_02746_),
    .B1(_02752_),
    .B2(_02759_),
    .Y(_03017_));
 sky130_fd_sc_hd__o2111ai_1 _27093_ (.A1(_06922_),
    .A2(_02748_),
    .B1(_02767_),
    .C1(_03011_),
    .D1(_03013_),
    .Y(_03018_));
 sky130_fd_sc_hd__a22o_1 _27094_ (.A1(_02753_),
    .A2(_02767_),
    .B1(_03011_),
    .B2(_03013_),
    .X(_03019_));
 sky130_fd_sc_hd__o211ai_2 _27095_ (.A1(net148),
    .A2(net147),
    .B1(_03018_),
    .C1(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__o2bb2ai_1 _27096_ (.A1_N(_03011_),
    .A2_N(_03013_),
    .B1(_03015_),
    .B2(_02755_),
    .Y(_03021_));
 sky130_fd_sc_hd__o211ai_2 _27097_ (.A1(_03004_),
    .A2(_03012_),
    .B1(_03011_),
    .C1(_03016_),
    .Y(_03022_));
 sky130_fd_sc_hd__o211ai_4 _27098_ (.A1(net148),
    .A2(net147),
    .B1(_03021_),
    .C1(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__o21ai_4 _27099_ (.A1(net146),
    .A2(_03010_),
    .B1(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__o31a_2 _27100_ (.A1(net148),
    .A2(net147),
    .A3(_03010_),
    .B1(_03023_),
    .X(_03026_));
 sky130_fd_sc_hd__and3_1 _27101_ (.A(_03024_),
    .B(_06921_),
    .C(_06919_),
    .X(_03027_));
 sky130_fd_sc_hd__o211ai_4 _27102_ (.A1(_03009_),
    .A2(net146),
    .B1(net226),
    .C1(_03020_),
    .Y(_03028_));
 sky130_fd_sc_hd__o221ai_4 _27103_ (.A1(_06918_),
    .A2(net249),
    .B1(net146),
    .B2(_03010_),
    .C1(_03023_),
    .Y(_03029_));
 sky130_fd_sc_hd__nand2_2 _27104_ (.A(_03028_),
    .B(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__nand4b_2 _27105_ (.A_N(_01850_),
    .B(_01852_),
    .C(_02162_),
    .D(_02165_),
    .Y(_03031_));
 sky130_fd_sc_hd__a21oi_1 _27106_ (.A1(_06315_),
    .A2(_02478_),
    .B1(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__nor3_1 _27107_ (.A(_02483_),
    .B(_03031_),
    .C(_02485_),
    .Y(_03033_));
 sky130_fd_sc_hd__o211ai_2 _27108_ (.A1(_06315_),
    .A2(_02478_),
    .B1(_03032_),
    .C1(_02775_),
    .Y(_03034_));
 sky130_fd_sc_hd__o211ai_4 _27109_ (.A1(_02780_),
    .A2(_02774_),
    .B1(_02776_),
    .C1(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__nand4_4 _27110_ (.A(_03033_),
    .B(_02776_),
    .C(_02775_),
    .D(_01862_),
    .Y(_03037_));
 sky130_fd_sc_hd__a21oi_2 _27111_ (.A1(_03035_),
    .A2(_03037_),
    .B1(_03030_),
    .Y(_03038_));
 sky130_fd_sc_hd__a21o_1 _27112_ (.A1(_03035_),
    .A2(_03037_),
    .B1(_03030_),
    .X(_03039_));
 sky130_fd_sc_hd__a31oi_2 _27113_ (.A1(_03030_),
    .A2(_03035_),
    .A3(_03037_),
    .B1(_09562_),
    .Y(_03040_));
 sky130_fd_sc_hd__a31o_1 _27114_ (.A1(_03030_),
    .A2(_03035_),
    .A3(_03037_),
    .B1(_09562_),
    .X(_03041_));
 sky130_fd_sc_hd__or3_1 _27115_ (.A(net156),
    .B(_09556_),
    .C(_03026_),
    .X(_03042_));
 sky130_fd_sc_hd__a22o_1 _27116_ (.A1(_03028_),
    .A2(_03029_),
    .B1(_03035_),
    .B2(_03037_),
    .X(_03043_));
 sky130_fd_sc_hd__o211ai_4 _27117_ (.A1(_03024_),
    .A2(net226),
    .B1(_03037_),
    .C1(_03035_),
    .Y(_03044_));
 sky130_fd_sc_hd__o221ai_4 _27118_ (.A1(net156),
    .A2(_09556_),
    .B1(_03027_),
    .B2(_03044_),
    .C1(_03043_),
    .Y(_03045_));
 sky130_fd_sc_hd__a2bb2oi_1 _27119_ (.A1_N(_09563_),
    .A2_N(_03024_),
    .B1(_03039_),
    .B2(_03040_),
    .Y(_03046_));
 sky130_fd_sc_hd__a22o_2 _27120_ (.A1(_09562_),
    .A2(_03026_),
    .B1(_03040_),
    .B2(_03039_),
    .X(_03048_));
 sky130_fd_sc_hd__o221a_2 _27121_ (.A1(_09563_),
    .A2(_03024_),
    .B1(_03038_),
    .B2(_03041_),
    .C1(_09578_),
    .X(_03049_));
 sky130_fd_sc_hd__a221o_1 _27122_ (.A1(_09562_),
    .A2(_03026_),
    .B1(_03040_),
    .B2(_03039_),
    .C1(net132),
    .X(_03050_));
 sky130_fd_sc_hd__nand3_4 _27123_ (.A(_03045_),
    .B(net235),
    .C(_03042_),
    .Y(_03051_));
 sky130_fd_sc_hd__o221a_1 _27124_ (.A1(_09563_),
    .A2(_03024_),
    .B1(_03038_),
    .B2(_03041_),
    .C1(net233),
    .X(_03052_));
 sky130_fd_sc_hd__o221ai_4 _27125_ (.A1(_09563_),
    .A2(_03024_),
    .B1(_03038_),
    .B2(_03041_),
    .C1(net233),
    .Y(_03053_));
 sky130_fd_sc_hd__o211ai_2 _27126_ (.A1(_06014_),
    .A2(_02495_),
    .B1(_02790_),
    .C1(_02794_),
    .Y(_03054_));
 sky130_fd_sc_hd__o21ai_4 _27127_ (.A1(_06314_),
    .A2(_02788_),
    .B1(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__a21oi_2 _27128_ (.A1(_03051_),
    .A2(_03053_),
    .B1(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__a21o_1 _27129_ (.A1(_03051_),
    .A2(_03053_),
    .B1(_03055_),
    .X(_03057_));
 sky130_fd_sc_hd__nand3_2 _27130_ (.A(_03051_),
    .B(_03053_),
    .C(_03055_),
    .Y(_03059_));
 sky130_fd_sc_hd__a31oi_2 _27131_ (.A1(_03051_),
    .A2(_03053_),
    .A3(_03055_),
    .B1(_09578_),
    .Y(_03060_));
 sky130_fd_sc_hd__a31o_1 _27132_ (.A1(_03051_),
    .A2(_03053_),
    .A3(_03055_),
    .B1(_09578_),
    .X(_03061_));
 sky130_fd_sc_hd__nand2_1 _27133_ (.A(_03060_),
    .B(_03057_),
    .Y(_03062_));
 sky130_fd_sc_hd__o22ai_4 _27134_ (.A1(net132),
    .A2(_03048_),
    .B1(_03056_),
    .B2(_03061_),
    .Y(_03063_));
 sky130_fd_sc_hd__o221a_1 _27135_ (.A1(_05767_),
    .A2(_02507_),
    .B1(_06013_),
    .B2(_02804_),
    .C1(_02525_),
    .X(_03064_));
 sky130_fd_sc_hd__o21ai_2 _27136_ (.A1(_02808_),
    .A2(_02812_),
    .B1(_02807_),
    .Y(_03065_));
 sky130_fd_sc_hd__a22o_1 _27137_ (.A1(_06311_),
    .A2(_06313_),
    .B1(_03060_),
    .B2(_03057_),
    .X(_03066_));
 sky130_fd_sc_hd__o221a_1 _27138_ (.A1(net132),
    .A2(_03048_),
    .B1(_03056_),
    .B2(_03061_),
    .C1(_06314_),
    .X(_03067_));
 sky130_fd_sc_hd__a211o_1 _27139_ (.A1(_03060_),
    .A2(_03057_),
    .B1(_03049_),
    .C1(_06315_),
    .X(_03068_));
 sky130_fd_sc_hd__a2bb2oi_2 _27140_ (.A1_N(net284),
    .A2_N(net281),
    .B1(_03050_),
    .B2(_03062_),
    .Y(_03070_));
 sky130_fd_sc_hd__o21ai_2 _27141_ (.A1(net284),
    .A2(net281),
    .B1(_03063_),
    .Y(_03071_));
 sky130_fd_sc_hd__o2111ai_1 _27142_ (.A1(_02812_),
    .A2(_02808_),
    .B1(_02807_),
    .C1(_03071_),
    .D1(_03068_),
    .Y(_03072_));
 sky130_fd_sc_hd__o21ai_1 _27143_ (.A1(_03067_),
    .A2(_03070_),
    .B1(_03065_),
    .Y(_03073_));
 sky130_fd_sc_hd__o211ai_1 _27144_ (.A1(_03049_),
    .A2(_03066_),
    .B1(_03071_),
    .C1(_03065_),
    .Y(_03074_));
 sky130_fd_sc_hd__o22ai_1 _27145_ (.A1(_02808_),
    .A2(_03064_),
    .B1(_03067_),
    .B2(_03070_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand3_2 _27146_ (.A(net131),
    .B(_03072_),
    .C(_03073_),
    .Y(_03076_));
 sky130_fd_sc_hd__a211o_1 _27147_ (.A1(_03050_),
    .A2(_03062_),
    .B1(net141),
    .C1(net140),
    .X(_03077_));
 sky130_fd_sc_hd__o211ai_1 _27148_ (.A1(net141),
    .A2(net140),
    .B1(_03074_),
    .C1(_03075_),
    .Y(_03078_));
 sky130_fd_sc_hd__o21ai_4 _27149_ (.A1(net131),
    .A2(_03063_),
    .B1(_03076_),
    .Y(_03079_));
 sky130_fd_sc_hd__and3_2 _27150_ (.A(_03078_),
    .B(_06013_),
    .C(_03077_),
    .X(_03081_));
 sky130_fd_sc_hd__o211ai_1 _27151_ (.A1(net285),
    .A2(_06012_),
    .B1(_03077_),
    .C1(_03078_),
    .Y(_03082_));
 sky130_fd_sc_hd__o211ai_4 _27152_ (.A1(net131),
    .A2(_03063_),
    .B1(_03076_),
    .C1(_06014_),
    .Y(_03083_));
 sky130_fd_sc_hd__o2bb2ai_1 _27153_ (.A1_N(_02820_),
    .A2_N(_02837_),
    .B1(_03079_),
    .B2(_06013_),
    .Y(_03084_));
 sky130_fd_sc_hd__a22oi_1 _27154_ (.A1(_02819_),
    .A2(_05768_),
    .B1(_03083_),
    .B2(_03082_),
    .Y(_03085_));
 sky130_fd_sc_hd__o21ai_1 _27155_ (.A1(_02821_),
    .A2(_02837_),
    .B1(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__o211ai_4 _27156_ (.A1(_03081_),
    .A2(_03084_),
    .B1(_03086_),
    .C1(_10954_),
    .Y(_03087_));
 sky130_fd_sc_hd__or3_1 _27157_ (.A(net137),
    .B(net135),
    .C(_03079_),
    .X(_03088_));
 sky130_fd_sc_hd__o31a_4 _27158_ (.A1(net137),
    .A2(net135),
    .A3(_03079_),
    .B1(_03087_),
    .X(_03089_));
 sky130_fd_sc_hd__or3_1 _27159_ (.A(_11459_),
    .B(net129),
    .C(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__a21oi_2 _27160_ (.A1(_03087_),
    .A2(_03088_),
    .B1(_05767_),
    .Y(_03092_));
 sky130_fd_sc_hd__o221a_1 _27161_ (.A1(_05765_),
    .A2(net288),
    .B1(_10954_),
    .B2(_03079_),
    .C1(_03087_),
    .X(_03093_));
 sky130_fd_sc_hd__o221ai_4 _27162_ (.A1(_05765_),
    .A2(net288),
    .B1(_10954_),
    .B2(_03079_),
    .C1(_03087_),
    .Y(_03094_));
 sky130_fd_sc_hd__nor2_1 _27163_ (.A(_03092_),
    .B(_03093_),
    .Y(_03095_));
 sky130_fd_sc_hd__and4_1 _27164_ (.A(_01909_),
    .B(_01911_),
    .C(_02244_),
    .D(_02245_),
    .X(_03096_));
 sky130_fd_sc_hd__nor3b_2 _27165_ (.A(_02544_),
    .B(_02546_),
    .C_N(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__nand3_1 _27166_ (.A(_02843_),
    .B(_03096_),
    .C(_02548_),
    .Y(_03098_));
 sky130_fd_sc_hd__o211a_1 _27167_ (.A1(_02846_),
    .A2(_02842_),
    .B1(_02844_),
    .C1(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__o211ai_2 _27168_ (.A1(_02846_),
    .A2(_02842_),
    .B1(_02844_),
    .C1(_03098_),
    .Y(_03100_));
 sky130_fd_sc_hd__nand4_2 _27169_ (.A(_03097_),
    .B(_02844_),
    .C(_02843_),
    .D(_01917_),
    .Y(_03101_));
 sky130_fd_sc_hd__a41oi_4 _27170_ (.A1(_01917_),
    .A2(_02843_),
    .A3(_02844_),
    .A4(_03097_),
    .B1(_03099_),
    .Y(_03103_));
 sky130_fd_sc_hd__nand2_1 _27171_ (.A(_03100_),
    .B(_03101_),
    .Y(_03104_));
 sky130_fd_sc_hd__o21ai_1 _27172_ (.A1(_03092_),
    .A2(_03093_),
    .B1(_03104_),
    .Y(_03105_));
 sky130_fd_sc_hd__nand2_1 _27173_ (.A(_03094_),
    .B(_03101_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand3_4 _27174_ (.A(_03094_),
    .B(_03100_),
    .C(_03101_),
    .Y(_03107_));
 sky130_fd_sc_hd__o221ai_4 _27175_ (.A1(_11459_),
    .A2(net129),
    .B1(_03092_),
    .B2(_03107_),
    .C1(_03105_),
    .Y(_03108_));
 sky130_fd_sc_hd__o311a_1 _27176_ (.A1(_11459_),
    .A2(net129),
    .A3(_03089_),
    .B1(_05507_),
    .C1(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__o2111ai_4 _27177_ (.A1(_03089_),
    .A2(_11465_),
    .B1(_05504_),
    .C1(_05502_),
    .D1(_03108_),
    .Y(_03110_));
 sky130_fd_sc_hd__a22o_1 _27178_ (.A1(_05502_),
    .A2(_05504_),
    .B1(_03090_),
    .B2(_03108_),
    .X(_03111_));
 sky130_fd_sc_hd__a21oi_1 _27179_ (.A1(_02854_),
    .A2(_02853_),
    .B1(_02851_),
    .Y(_03112_));
 sky130_fd_sc_hd__a221oi_2 _27180_ (.A1(_02854_),
    .A2(_02853_),
    .B1(_03111_),
    .B2(_03110_),
    .C1(_02851_),
    .Y(_03114_));
 sky130_fd_sc_hd__o221ai_4 _27181_ (.A1(_11465_),
    .A2(_03089_),
    .B1(_11944_),
    .B2(_03114_),
    .C1(_03108_),
    .Y(_03115_));
 sky130_fd_sc_hd__a21oi_1 _27182_ (.A1(_05119_),
    .A2(_02859_),
    .B1(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__o311a_1 _27183_ (.A1(_02260_),
    .A2(_02559_),
    .A3(_02856_),
    .B1(_03115_),
    .C1(_05119_),
    .X(_03117_));
 sky130_fd_sc_hd__nor2_1 _27184_ (.A(_03116_),
    .B(_03117_),
    .Y(net105));
 sky130_fd_sc_hd__o21ai_1 _27185_ (.A1(_02859_),
    .A2(_03115_),
    .B1(_05119_),
    .Y(_03118_));
 sky130_fd_sc_hd__and4_1 _27186_ (.A(_02106_),
    .B(_02107_),
    .C(_02418_),
    .D(_02420_),
    .X(_03119_));
 sky130_fd_sc_hd__nand3_1 _27187_ (.A(_02982_),
    .B(_03119_),
    .C(_02723_),
    .Y(_03120_));
 sky130_fd_sc_hd__o211ai_4 _27188_ (.A1(_02986_),
    .A2(_02980_),
    .B1(_02984_),
    .C1(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__and4_1 _27189_ (.A(_03119_),
    .B(_02722_),
    .C(_02720_),
    .D(_02116_),
    .X(_03122_));
 sky130_fd_sc_hd__nand3_4 _27190_ (.A(_03122_),
    .B(_02984_),
    .C(_02982_),
    .Y(_03124_));
 sky130_fd_sc_hd__nand2_1 _27191_ (.A(_03121_),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__o211ai_4 _27192_ (.A1(_02867_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_02875_),
    .Y(_03126_));
 sky130_fd_sc_hd__o21ai_2 _27193_ (.A1(net260),
    .A2(net255),
    .B1(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__or3_1 _27194_ (.A(net239),
    .B(_06292_),
    .C(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__and3_1 _27195_ (.A(net240),
    .B(_10971_),
    .C(_03126_),
    .X(_03129_));
 sky130_fd_sc_hd__a21o_1 _27196_ (.A1(_10963_),
    .A2(_10964_),
    .B1(_03127_),
    .X(_03130_));
 sky130_fd_sc_hd__and3_1 _27197_ (.A(_10963_),
    .B(_10964_),
    .C(_03127_),
    .X(_03131_));
 sky130_fd_sc_hd__a22o_1 _27198_ (.A1(_10966_),
    .A2(_10968_),
    .B1(_03126_),
    .B2(net240),
    .X(_03132_));
 sky130_fd_sc_hd__o211ai_2 _27199_ (.A1(_02887_),
    .A2(_02612_),
    .B1(_02604_),
    .C1(_02880_),
    .Y(_03133_));
 sky130_fd_sc_hd__o2111ai_4 _27200_ (.A1(_10492_),
    .A2(_02878_),
    .B1(_03130_),
    .C1(_03132_),
    .D1(_03133_),
    .Y(_03135_));
 sky130_fd_sc_hd__o221ai_4 _27201_ (.A1(_03129_),
    .A2(_03131_),
    .B1(_02881_),
    .B2(_02888_),
    .C1(_02880_),
    .Y(_03136_));
 sky130_fd_sc_hd__o211ai_2 _27202_ (.A1(net239),
    .A2(_06292_),
    .B1(_03135_),
    .C1(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__a21oi_1 _27203_ (.A1(net240),
    .A2(_03126_),
    .B1(_06293_),
    .Y(_03138_));
 sky130_fd_sc_hd__a2bb2oi_1 _27204_ (.A1_N(net239),
    .A2_N(_06292_),
    .B1(_03135_),
    .B2(_03136_),
    .Y(_03139_));
 sky130_fd_sc_hd__o21a_2 _27205_ (.A1(_06293_),
    .A2(_03127_),
    .B1(_03137_),
    .X(_03140_));
 sky130_fd_sc_hd__a2bb2oi_1 _27206_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_03128_),
    .B2(_03137_),
    .Y(_03141_));
 sky130_fd_sc_hd__a31oi_2 _27207_ (.A1(_03136_),
    .A2(_06293_),
    .A3(_03135_),
    .B1(_10492_),
    .Y(_03142_));
 sky130_fd_sc_hd__o21ai_1 _27208_ (.A1(_06293_),
    .A2(_03127_),
    .B1(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__a21oi_2 _27209_ (.A1(_03128_),
    .A2(_03142_),
    .B1(_03141_),
    .Y(_03144_));
 sky130_fd_sc_hd__o41ai_2 _27210_ (.A1(net164),
    .A2(_10490_),
    .A3(_03138_),
    .A4(_03139_),
    .B1(_03143_),
    .Y(_03146_));
 sky130_fd_sc_hd__o21ai_1 _27211_ (.A1(net151),
    .A2(_02895_),
    .B1(_02908_),
    .Y(_03147_));
 sky130_fd_sc_hd__o211ai_2 _27212_ (.A1(_02895_),
    .A2(net151),
    .B1(_02908_),
    .C1(_02906_),
    .Y(_03148_));
 sky130_fd_sc_hd__o22ai_2 _27213_ (.A1(net152),
    .A2(_02896_),
    .B1(_03147_),
    .B2(_02905_),
    .Y(_03149_));
 sky130_fd_sc_hd__a21oi_4 _27214_ (.A1(_02897_),
    .A2(_03148_),
    .B1(_03146_),
    .Y(_03150_));
 sky130_fd_sc_hd__nand2_1 _27215_ (.A(_03144_),
    .B(_03149_),
    .Y(_03151_));
 sky130_fd_sc_hd__a21oi_1 _27216_ (.A1(_03128_),
    .A2(_03137_),
    .B1(net209),
    .Y(_03152_));
 sky130_fd_sc_hd__o22ai_4 _27217_ (.A1(net238),
    .A2(net236),
    .B1(_03144_),
    .B2(_03149_),
    .Y(_03153_));
 sky130_fd_sc_hd__o22ai_2 _27218_ (.A1(net209),
    .A2(_03140_),
    .B1(_03150_),
    .B2(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__o22a_1 _27219_ (.A1(net209),
    .A2(_03140_),
    .B1(_03150_),
    .B2(_03153_),
    .X(_03155_));
 sky130_fd_sc_hd__and3_2 _27220_ (.A(_03154_),
    .B(_06902_),
    .C(_06900_),
    .X(_03157_));
 sky130_fd_sc_hd__or3_1 _27221_ (.A(net229),
    .B(net228),
    .C(_03155_),
    .X(_03158_));
 sky130_fd_sc_hd__and3_1 _27222_ (.A(_02037_),
    .B(_02352_),
    .C(_02354_),
    .X(_03159_));
 sky130_fd_sc_hd__nand4_1 _27223_ (.A(_02034_),
    .B(_02036_),
    .C(_02352_),
    .D(_02354_),
    .Y(_03160_));
 sky130_fd_sc_hd__a211oi_1 _27224_ (.A1(_02626_),
    .A2(_02647_),
    .B1(_03160_),
    .C1(_02651_),
    .Y(_03161_));
 sky130_fd_sc_hd__nand2_1 _27225_ (.A(_02922_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__o211a_1 _27226_ (.A1(_02925_),
    .A2(_02921_),
    .B1(_02923_),
    .C1(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__o211ai_4 _27227_ (.A1(_02925_),
    .A2(_02921_),
    .B1(_02923_),
    .C1(_03162_),
    .Y(_03164_));
 sky130_fd_sc_hd__o2111a_1 _27228_ (.A1(_02044_),
    .A2(_02047_),
    .B1(_02650_),
    .C1(_03159_),
    .D1(_02653_),
    .X(_03165_));
 sky130_fd_sc_hd__nand3_4 _27229_ (.A(_03165_),
    .B(_02923_),
    .C(_02922_),
    .Y(_03166_));
 sky130_fd_sc_hd__o21a_1 _27230_ (.A1(net170),
    .A2(net168),
    .B1(_03154_),
    .X(_03168_));
 sky130_fd_sc_hd__o21ai_2 _27231_ (.A1(net170),
    .A2(net168),
    .B1(_03154_),
    .Y(_03169_));
 sky130_fd_sc_hd__o22ai_1 _27232_ (.A1(net167),
    .A2(_10024_),
    .B1(_03150_),
    .B2(_03153_),
    .Y(_03170_));
 sky130_fd_sc_hd__o221a_1 _27233_ (.A1(net209),
    .A2(_03140_),
    .B1(_03150_),
    .B2(_03153_),
    .C1(net152),
    .X(_03171_));
 sky130_fd_sc_hd__o221ai_4 _27234_ (.A1(net209),
    .A2(_03140_),
    .B1(_03150_),
    .B2(_03153_),
    .C1(net152),
    .Y(_03172_));
 sky130_fd_sc_hd__a22oi_2 _27235_ (.A1(_03164_),
    .A2(_03166_),
    .B1(_03169_),
    .B2(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__o2bb2ai_4 _27236_ (.A1_N(_03164_),
    .A2_N(_03166_),
    .B1(_03168_),
    .B2(_03171_),
    .Y(_03174_));
 sky130_fd_sc_hd__o211ai_1 _27237_ (.A1(_03170_),
    .A2(_03152_),
    .B1(_03166_),
    .C1(_03169_),
    .Y(_03175_));
 sky130_fd_sc_hd__nand4_4 _27238_ (.A(_03164_),
    .B(_03166_),
    .C(_03169_),
    .D(_03172_),
    .Y(_03176_));
 sky130_fd_sc_hd__o22ai_2 _27239_ (.A1(net229),
    .A2(net228),
    .B1(_03175_),
    .B2(_03163_),
    .Y(_03177_));
 sky130_fd_sc_hd__nand3_1 _27240_ (.A(_03174_),
    .B(_03176_),
    .C(_06903_),
    .Y(_03180_));
 sky130_fd_sc_hd__a31oi_4 _27241_ (.A1(_03174_),
    .A2(_03176_),
    .A3(_06903_),
    .B1(_03157_),
    .Y(_03181_));
 sky130_fd_sc_hd__o22ai_4 _27242_ (.A1(_06903_),
    .A2(_03155_),
    .B1(_03173_),
    .B2(_03177_),
    .Y(_03182_));
 sky130_fd_sc_hd__and3_1 _27243_ (.A(_07228_),
    .B(_07230_),
    .C(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__or3_1 _27244_ (.A(net207),
    .B(net204),
    .C(_03181_),
    .X(_03184_));
 sky130_fd_sc_hd__a311oi_4 _27245_ (.A1(_03174_),
    .A2(_03176_),
    .A3(_06903_),
    .B1(net171),
    .C1(_03157_),
    .Y(_03185_));
 sky130_fd_sc_hd__nand3_2 _27246_ (.A(_03180_),
    .B(_09594_),
    .C(_03158_),
    .Y(_03186_));
 sky130_fd_sc_hd__a2bb2oi_1 _27247_ (.A1_N(net189),
    .A2_N(net188),
    .B1(_03158_),
    .B2(_03180_),
    .Y(_03187_));
 sky130_fd_sc_hd__o21ai_4 _27248_ (.A1(net189),
    .A2(net188),
    .B1(_03182_),
    .Y(_03188_));
 sky130_fd_sc_hd__o21ai_1 _27249_ (.A1(_02935_),
    .A2(_02934_),
    .B1(_02939_),
    .Y(_03189_));
 sky130_fd_sc_hd__a21oi_2 _27250_ (.A1(_02933_),
    .A2(_02936_),
    .B1(_02938_),
    .Y(_03191_));
 sky130_fd_sc_hd__o21a_1 _27251_ (.A1(_03185_),
    .A2(_03187_),
    .B1(_03191_),
    .X(_03192_));
 sky130_fd_sc_hd__o21ai_2 _27252_ (.A1(_03185_),
    .A2(_03187_),
    .B1(_03191_),
    .Y(_03193_));
 sky130_fd_sc_hd__o21ai_1 _27253_ (.A1(_09594_),
    .A2(_03181_),
    .B1(_03189_),
    .Y(_03194_));
 sky130_fd_sc_hd__nand3_1 _27254_ (.A(_03186_),
    .B(_03188_),
    .C(_03189_),
    .Y(_03195_));
 sky130_fd_sc_hd__o22ai_2 _27255_ (.A1(net207),
    .A2(net204),
    .B1(_03185_),
    .B2(_03194_),
    .Y(_03196_));
 sky130_fd_sc_hd__o211ai_2 _27256_ (.A1(_03194_),
    .A2(_03185_),
    .B1(_07233_),
    .C1(_03193_),
    .Y(_03197_));
 sky130_fd_sc_hd__o22ai_4 _27257_ (.A1(_07233_),
    .A2(_03181_),
    .B1(_03192_),
    .B2(_03196_),
    .Y(_03198_));
 sky130_fd_sc_hd__o211a_1 _27258_ (.A1(_02677_),
    .A2(net201),
    .B1(_02952_),
    .C1(_02693_),
    .X(_03199_));
 sky130_fd_sc_hd__o221ai_1 _27259_ (.A1(net201),
    .A2(_02677_),
    .B1(net178),
    .B2(_02949_),
    .C1(_02693_),
    .Y(_03200_));
 sky130_fd_sc_hd__o2bb2ai_1 _27260_ (.A1_N(_02679_),
    .A2_N(_02693_),
    .B1(_02947_),
    .B2(_08731_),
    .Y(_03202_));
 sky130_fd_sc_hd__a31oi_2 _27261_ (.A1(_02679_),
    .A2(_02693_),
    .A3(_02952_),
    .B1(_02953_),
    .Y(_03203_));
 sky130_fd_sc_hd__a31o_1 _27262_ (.A1(_07233_),
    .A2(_03193_),
    .A3(_03195_),
    .B1(_09140_),
    .X(_03204_));
 sky130_fd_sc_hd__a311oi_2 _27263_ (.A1(_07233_),
    .A2(_03193_),
    .A3(_03195_),
    .B1(_09140_),
    .C1(_03183_),
    .Y(_03205_));
 sky130_fd_sc_hd__nand3_1 _27264_ (.A(_03197_),
    .B(_09139_),
    .C(_03184_),
    .Y(_03206_));
 sky130_fd_sc_hd__a2bb2oi_2 _27265_ (.A1_N(net194),
    .A2_N(net191),
    .B1(_03184_),
    .B2(_03197_),
    .Y(_03207_));
 sky130_fd_sc_hd__o21ai_1 _27266_ (.A1(net194),
    .A2(net191),
    .B1(_03198_),
    .Y(_03208_));
 sky130_fd_sc_hd__nor2_1 _27267_ (.A(_03205_),
    .B(_03207_),
    .Y(_03209_));
 sky130_fd_sc_hd__o2111ai_1 _27268_ (.A1(net178),
    .A2(_02949_),
    .B1(_03202_),
    .C1(_03206_),
    .D1(_03208_),
    .Y(_03210_));
 sky130_fd_sc_hd__o2bb2ai_1 _27269_ (.A1_N(_02952_),
    .A2_N(_03202_),
    .B1(_03205_),
    .B2(_03207_),
    .Y(_03211_));
 sky130_fd_sc_hd__nand3_2 _27270_ (.A(_03211_),
    .B(_07548_),
    .C(_03210_),
    .Y(_03213_));
 sky130_fd_sc_hd__a211o_1 _27271_ (.A1(_03184_),
    .A2(_03197_),
    .B1(_07544_),
    .C1(_07546_),
    .X(_03214_));
 sky130_fd_sc_hd__o211ai_1 _27272_ (.A1(_03183_),
    .A2(_03204_),
    .B1(_03203_),
    .C1(_03208_),
    .Y(_03215_));
 sky130_fd_sc_hd__o22ai_1 _27273_ (.A1(_02953_),
    .A2(_03199_),
    .B1(_03205_),
    .B2(_03207_),
    .Y(_03216_));
 sky130_fd_sc_hd__nand3_1 _27274_ (.A(_03216_),
    .B(_07548_),
    .C(_03215_),
    .Y(_03217_));
 sky130_fd_sc_hd__o21a_1 _27275_ (.A1(_07548_),
    .A2(_03198_),
    .B1(_03213_),
    .X(_03218_));
 sky130_fd_sc_hd__o21ai_4 _27276_ (.A1(_07548_),
    .A2(_03198_),
    .B1(_03213_),
    .Y(_03219_));
 sky130_fd_sc_hd__o211ai_4 _27277_ (.A1(_03198_),
    .A2(_07548_),
    .B1(_08731_),
    .C1(_03213_),
    .Y(_03220_));
 sky130_fd_sc_hd__and3_1 _27278_ (.A(_03217_),
    .B(net178),
    .C(_03214_),
    .X(_03221_));
 sky130_fd_sc_hd__nand3_2 _27279_ (.A(_03217_),
    .B(net178),
    .C(_03214_),
    .Y(_03222_));
 sky130_fd_sc_hd__nand2_1 _27280_ (.A(_03220_),
    .B(_03222_),
    .Y(_03224_));
 sky130_fd_sc_hd__o2bb2ai_1 _27281_ (.A1_N(_02864_),
    .A2_N(_02865_),
    .B1(_02965_),
    .B2(net201),
    .Y(_03225_));
 sky130_fd_sc_hd__nand3_2 _27282_ (.A(_02864_),
    .B(_02865_),
    .C(_02969_),
    .Y(_03226_));
 sky130_fd_sc_hd__a31oi_2 _27283_ (.A1(_02864_),
    .A2(_02865_),
    .A3(_02969_),
    .B1(_02966_),
    .Y(_03227_));
 sky130_fd_sc_hd__o2111ai_1 _27284_ (.A1(net201),
    .A2(_02965_),
    .B1(_03220_),
    .C1(_03222_),
    .D1(_03226_),
    .Y(_03228_));
 sky130_fd_sc_hd__a22o_1 _27285_ (.A1(_03220_),
    .A2(_03222_),
    .B1(_03226_),
    .B2(_02967_),
    .X(_03229_));
 sky130_fd_sc_hd__nand3_2 _27286_ (.A(_03229_),
    .B(_07916_),
    .C(_03228_),
    .Y(_03230_));
 sky130_fd_sc_hd__o211ai_1 _27287_ (.A1(_02965_),
    .A2(net201),
    .B1(_03226_),
    .C1(_03224_),
    .Y(_03231_));
 sky130_fd_sc_hd__o2111ai_4 _27288_ (.A1(net197),
    .A2(_02964_),
    .B1(_03220_),
    .C1(_03222_),
    .D1(_03225_),
    .Y(_03232_));
 sky130_fd_sc_hd__a21oi_1 _27289_ (.A1(_03224_),
    .A2(_03227_),
    .B1(_07917_),
    .Y(_03233_));
 sky130_fd_sc_hd__o211ai_2 _27290_ (.A1(net183),
    .A2(net182),
    .B1(_03231_),
    .C1(_03232_),
    .Y(_03235_));
 sky130_fd_sc_hd__o2bb2a_4 _27291_ (.A1_N(_03233_),
    .A2_N(_03232_),
    .B1(_03219_),
    .B2(_07916_),
    .X(_03236_));
 sky130_fd_sc_hd__o211a_1 _27292_ (.A1(_07916_),
    .A2(_03218_),
    .B1(_03230_),
    .C1(net197),
    .X(_03237_));
 sky130_fd_sc_hd__o211ai_4 _27293_ (.A1(_07916_),
    .A2(_03218_),
    .B1(_03230_),
    .C1(net197),
    .Y(_03238_));
 sky130_fd_sc_hd__o211a_1 _27294_ (.A1(net162),
    .A2(_03219_),
    .B1(net201),
    .C1(_03235_),
    .X(_03239_));
 sky130_fd_sc_hd__o211ai_4 _27295_ (.A1(net162),
    .A2(_03219_),
    .B1(net201),
    .C1(_03235_),
    .Y(_03240_));
 sky130_fd_sc_hd__nand2_1 _27296_ (.A(_03238_),
    .B(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand3_1 _27297_ (.A(_03121_),
    .B(_03124_),
    .C(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__a21o_1 _27298_ (.A1(_03121_),
    .A2(_03124_),
    .B1(_03241_),
    .X(_03243_));
 sky130_fd_sc_hd__o2bb2ai_1 _27299_ (.A1_N(_03121_),
    .A2_N(_03124_),
    .B1(_03237_),
    .B2(_03239_),
    .Y(_03244_));
 sky130_fd_sc_hd__nand4_1 _27300_ (.A(_03121_),
    .B(_03124_),
    .C(_03238_),
    .D(_03240_),
    .Y(_03246_));
 sky130_fd_sc_hd__nand3_4 _27301_ (.A(_03244_),
    .B(_03246_),
    .C(net159),
    .Y(_03247_));
 sky130_fd_sc_hd__or3_1 _27302_ (.A(net181),
    .B(net179),
    .C(_03236_),
    .X(_03248_));
 sky130_fd_sc_hd__a221o_1 _27303_ (.A1(_07917_),
    .A2(_03218_),
    .B1(_03233_),
    .B2(_03232_),
    .C1(net159),
    .X(_03249_));
 sky130_fd_sc_hd__nand3_1 _27304_ (.A(_03243_),
    .B(net159),
    .C(_03242_),
    .Y(_03250_));
 sky130_fd_sc_hd__o21ai_1 _27305_ (.A1(net159),
    .A2(_03236_),
    .B1(_03247_),
    .Y(_03251_));
 sky130_fd_sc_hd__and3_1 _27306_ (.A(_08715_),
    .B(_03249_),
    .C(_03250_),
    .X(_03252_));
 sky130_fd_sc_hd__a22o_2 _27307_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_03247_),
    .B2(_03248_),
    .X(_03253_));
 sky130_fd_sc_hd__o311a_1 _27308_ (.A1(net181),
    .A2(net179),
    .A3(_03236_),
    .B1(_07935_),
    .C1(_03247_),
    .X(_03254_));
 sky130_fd_sc_hd__o211ai_4 _27309_ (.A1(net159),
    .A2(_03236_),
    .B1(_07935_),
    .C1(_03247_),
    .Y(_03255_));
 sky130_fd_sc_hd__o211ai_4 _27310_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_03249_),
    .C1(_03250_),
    .Y(_03257_));
 sky130_fd_sc_hd__a21oi_1 _27311_ (.A1(_02736_),
    .A2(_02993_),
    .B1(_02998_),
    .Y(_03258_));
 sky130_fd_sc_hd__o211a_1 _27312_ (.A1(net223),
    .A2(_02732_),
    .B1(_02993_),
    .C1(_02997_),
    .X(_03259_));
 sky130_fd_sc_hd__a31o_1 _27313_ (.A1(_02736_),
    .A2(_02993_),
    .A3(_02997_),
    .B1(_02998_),
    .X(_03260_));
 sky130_fd_sc_hd__a31oi_2 _27314_ (.A1(_02736_),
    .A2(_02993_),
    .A3(_02997_),
    .B1(_02998_),
    .Y(_03261_));
 sky130_fd_sc_hd__a21oi_1 _27315_ (.A1(_03255_),
    .A2(_03257_),
    .B1(_03260_),
    .Y(_03262_));
 sky130_fd_sc_hd__o2bb2ai_4 _27316_ (.A1_N(_03255_),
    .A2_N(_03257_),
    .B1(_03258_),
    .B2(_02996_),
    .Y(_03263_));
 sky130_fd_sc_hd__o211a_1 _27317_ (.A1(_02998_),
    .A2(_03259_),
    .B1(_03257_),
    .C1(_03255_),
    .X(_03264_));
 sky130_fd_sc_hd__o211ai_4 _27318_ (.A1(_02998_),
    .A2(_03259_),
    .B1(_03257_),
    .C1(_03255_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand3_1 _27319_ (.A(_03263_),
    .B(_03265_),
    .C(net149),
    .Y(_03266_));
 sky130_fd_sc_hd__o311a_1 _27320_ (.A1(net181),
    .A2(_03236_),
    .A3(net179),
    .B1(_08715_),
    .C1(_03247_),
    .X(_03268_));
 sky130_fd_sc_hd__a21oi_1 _27321_ (.A1(_03263_),
    .A2(_03265_),
    .B1(_08715_),
    .Y(_03269_));
 sky130_fd_sc_hd__o22ai_1 _27322_ (.A1(net157),
    .A2(_08712_),
    .B1(_03262_),
    .B2(_03264_),
    .Y(_03270_));
 sky130_fd_sc_hd__a31o_1 _27323_ (.A1(_08715_),
    .A2(_03247_),
    .A3(_03248_),
    .B1(_03269_),
    .X(_03271_));
 sky130_fd_sc_hd__inv_2 _27324_ (.A(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__o21ai_2 _27325_ (.A1(_07246_),
    .A2(_03010_),
    .B1(_03017_),
    .Y(_03273_));
 sky130_fd_sc_hd__a2bb2oi_1 _27326_ (.A1_N(_03012_),
    .A2_N(_03004_),
    .B1(_03011_),
    .B2(_03017_),
    .Y(_03274_));
 sky130_fd_sc_hd__a31oi_2 _27327_ (.A1(_03263_),
    .A2(_03265_),
    .A3(net149),
    .B1(_07565_),
    .Y(_03275_));
 sky130_fd_sc_hd__a311oi_4 _27328_ (.A1(_03263_),
    .A2(_03265_),
    .A3(net149),
    .B1(_03252_),
    .C1(_07565_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand3_1 _27329_ (.A(_03266_),
    .B(_07564_),
    .C(_03253_),
    .Y(_03277_));
 sky130_fd_sc_hd__a2bb2oi_4 _27330_ (.A1_N(net221),
    .A2_N(net219),
    .B1(_03253_),
    .B2(_03266_),
    .Y(_03279_));
 sky130_fd_sc_hd__o221ai_2 _27331_ (.A1(net221),
    .A2(net219),
    .B1(net149),
    .B2(_03251_),
    .C1(_03270_),
    .Y(_03280_));
 sky130_fd_sc_hd__a211oi_2 _27332_ (.A1(_03013_),
    .A2(_03273_),
    .B1(_03276_),
    .C1(_03279_),
    .Y(_03281_));
 sky130_fd_sc_hd__o21ai_1 _27333_ (.A1(_03276_),
    .A2(_03279_),
    .B1(_03274_),
    .Y(_03282_));
 sky130_fd_sc_hd__o21ai_2 _27334_ (.A1(net148),
    .A2(net147),
    .B1(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__nand3_1 _27335_ (.A(_03280_),
    .B(_03274_),
    .C(_03277_),
    .Y(_03284_));
 sky130_fd_sc_hd__o2bb2ai_1 _27336_ (.A1_N(_03013_),
    .A2_N(_03273_),
    .B1(_03276_),
    .B2(_03279_),
    .Y(_03285_));
 sky130_fd_sc_hd__or4_1 _27337_ (.A(net148),
    .B(net147),
    .C(_03268_),
    .D(_03269_),
    .X(_03286_));
 sky130_fd_sc_hd__o211ai_4 _27338_ (.A1(net148),
    .A2(net147),
    .B1(_03284_),
    .C1(_03285_),
    .Y(_03287_));
 sky130_fd_sc_hd__o22a_2 _27339_ (.A1(net146),
    .A2(_03272_),
    .B1(_03281_),
    .B2(_03283_),
    .X(_03288_));
 sky130_fd_sc_hd__o311a_1 _27340_ (.A1(net145),
    .A2(_03268_),
    .A3(_03269_),
    .B1(_07246_),
    .C1(_03287_),
    .X(_03291_));
 sky130_fd_sc_hd__o211ai_4 _27341_ (.A1(net146),
    .A2(_03271_),
    .B1(_07246_),
    .C1(_03287_),
    .Y(_03292_));
 sky130_fd_sc_hd__a21oi_1 _27342_ (.A1(_03286_),
    .A2(_03287_),
    .B1(_07246_),
    .Y(_03293_));
 sky130_fd_sc_hd__o221ai_4 _27343_ (.A1(net146),
    .A2(_03272_),
    .B1(_03281_),
    .B2(_03283_),
    .C1(net223),
    .Y(_03294_));
 sky130_fd_sc_hd__o2111a_1 _27344_ (.A1(_03026_),
    .A2(_06922_),
    .B1(_03292_),
    .C1(_03044_),
    .D1(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__o2111ai_4 _27345_ (.A1(_03026_),
    .A2(_06922_),
    .B1(_03292_),
    .C1(_03044_),
    .D1(_03294_),
    .Y(_03296_));
 sky130_fd_sc_hd__a22oi_1 _27346_ (.A1(_03028_),
    .A2(_03044_),
    .B1(_03292_),
    .B2(_03294_),
    .Y(_03297_));
 sky130_fd_sc_hd__o2bb2ai_2 _27347_ (.A1_N(_03028_),
    .A2_N(_03044_),
    .B1(_03291_),
    .B2(_03293_),
    .Y(_03298_));
 sky130_fd_sc_hd__o2111ai_2 _27348_ (.A1(_09551_),
    .A2(_09558_),
    .B1(_09561_),
    .C1(_03296_),
    .D1(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__o221a_2 _27349_ (.A1(net146),
    .A2(_03272_),
    .B1(_03281_),
    .B2(_03283_),
    .C1(_09562_),
    .X(_03300_));
 sky130_fd_sc_hd__inv_2 _27350_ (.A(_03300_),
    .Y(_03302_));
 sky130_fd_sc_hd__a2bb2oi_2 _27351_ (.A1_N(net156),
    .A2_N(_09556_),
    .B1(_03296_),
    .B2(_03298_),
    .Y(_03303_));
 sky130_fd_sc_hd__o22ai_2 _27352_ (.A1(net156),
    .A2(net154),
    .B1(_03295_),
    .B2(_03297_),
    .Y(_03304_));
 sky130_fd_sc_hd__o21ai_2 _27353_ (.A1(net144),
    .A2(_03288_),
    .B1(_03299_),
    .Y(_03305_));
 sky130_fd_sc_hd__o211a_2 _27354_ (.A1(_03288_),
    .A2(net144),
    .B1(net226),
    .C1(_03299_),
    .X(_03306_));
 sky130_fd_sc_hd__o21ai_4 _27355_ (.A1(_03300_),
    .A2(_03303_),
    .B1(net226),
    .Y(_03307_));
 sky130_fd_sc_hd__o211ai_4 _27356_ (.A1(_06918_),
    .A2(net249),
    .B1(_03302_),
    .C1(_03304_),
    .Y(_03308_));
 sky130_fd_sc_hd__o211a_1 _27357_ (.A1(_02184_),
    .A2(_02175_),
    .B1(_02183_),
    .C1(_02498_),
    .X(_03309_));
 sky130_fd_sc_hd__o2111a_1 _27358_ (.A1(_06014_),
    .A2(_02495_),
    .B1(_02794_),
    .C1(_03309_),
    .D1(_02797_),
    .X(_03310_));
 sky130_fd_sc_hd__nand4_1 _27359_ (.A(_02797_),
    .B(_02502_),
    .C(_02187_),
    .D(_02794_),
    .Y(_03311_));
 sky130_fd_sc_hd__a31oi_1 _27360_ (.A1(_03045_),
    .A2(net235),
    .A3(_03042_),
    .B1(_03311_),
    .Y(_03313_));
 sky130_fd_sc_hd__o21ai_1 _27361_ (.A1(net233),
    .A2(_03046_),
    .B1(_03310_),
    .Y(_03314_));
 sky130_fd_sc_hd__a21oi_1 _27362_ (.A1(_03051_),
    .A2(_03310_),
    .B1(_03052_),
    .Y(_03315_));
 sky130_fd_sc_hd__a211oi_1 _27363_ (.A1(_03055_),
    .A2(_03051_),
    .B1(_03052_),
    .C1(_03313_),
    .Y(_03316_));
 sky130_fd_sc_hd__o211ai_4 _27364_ (.A1(_03048_),
    .A2(net235),
    .B1(_03314_),
    .C1(_03059_),
    .Y(_03317_));
 sky130_fd_sc_hd__o2111a_1 _27365_ (.A1(_02771_),
    .A2(_02792_),
    .B1(_02202_),
    .C1(_02502_),
    .D1(_02797_),
    .X(_03318_));
 sky130_fd_sc_hd__nand3_4 _27366_ (.A(_03051_),
    .B(_03318_),
    .C(_03053_),
    .Y(_03319_));
 sky130_fd_sc_hd__a31o_1 _27367_ (.A1(_03051_),
    .A2(_03053_),
    .A3(_03318_),
    .B1(_03316_),
    .X(_03320_));
 sky130_fd_sc_hd__a22oi_4 _27368_ (.A1(_03307_),
    .A2(_03308_),
    .B1(_03317_),
    .B2(_03319_),
    .Y(_03321_));
 sky130_fd_sc_hd__a22o_1 _27369_ (.A1(_03307_),
    .A2(_03308_),
    .B1(_03317_),
    .B2(_03319_),
    .X(_03322_));
 sky130_fd_sc_hd__o31a_1 _27370_ (.A1(net226),
    .A2(_03300_),
    .A3(_03303_),
    .B1(_03319_),
    .X(_03324_));
 sky130_fd_sc_hd__o31ai_2 _27371_ (.A1(net226),
    .A2(_03300_),
    .A3(_03303_),
    .B1(_03319_),
    .Y(_03325_));
 sky130_fd_sc_hd__nand3_2 _27372_ (.A(_03308_),
    .B(_03317_),
    .C(_03319_),
    .Y(_03326_));
 sky130_fd_sc_hd__a211oi_4 _27373_ (.A1(_03315_),
    .A2(_03059_),
    .B1(_03306_),
    .C1(_03325_),
    .Y(_03327_));
 sky130_fd_sc_hd__o221ai_4 _27374_ (.A1(net142),
    .A2(_09573_),
    .B1(_03306_),
    .B2(_03326_),
    .C1(_03322_),
    .Y(_03328_));
 sky130_fd_sc_hd__or3_4 _27375_ (.A(net142),
    .B(_09573_),
    .C(_03305_),
    .X(_03329_));
 sky130_fd_sc_hd__o31a_4 _27376_ (.A1(_09578_),
    .A2(_03321_),
    .A3(_03327_),
    .B1(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__o31ai_4 _27377_ (.A1(_09578_),
    .A2(_03321_),
    .A3(_03327_),
    .B1(_03329_),
    .Y(_03331_));
 sky130_fd_sc_hd__or3_1 _27378_ (.A(net141),
    .B(net140),
    .C(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__o211a_1 _27379_ (.A1(_02812_),
    .A2(_02808_),
    .B1(_02807_),
    .C1(_03071_),
    .X(_03333_));
 sky130_fd_sc_hd__o22a_1 _27380_ (.A1(_03049_),
    .A2(_03066_),
    .B1(_03070_),
    .B2(_03065_),
    .X(_03335_));
 sky130_fd_sc_hd__a21oi_2 _27381_ (.A1(_03065_),
    .A2(_03068_),
    .B1(_03070_),
    .Y(_03336_));
 sky130_fd_sc_hd__o31a_1 _27382_ (.A1(_09578_),
    .A2(_03321_),
    .A3(_03327_),
    .B1(_06629_),
    .X(_03337_));
 sky130_fd_sc_hd__o311a_2 _27383_ (.A1(_09578_),
    .A2(_03321_),
    .A3(_03327_),
    .B1(_03329_),
    .C1(_06629_),
    .X(_03338_));
 sky130_fd_sc_hd__nand3_1 _27384_ (.A(_03328_),
    .B(_03329_),
    .C(_06629_),
    .Y(_03339_));
 sky130_fd_sc_hd__a22oi_4 _27385_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_03328_),
    .B2(_03329_),
    .Y(_03340_));
 sky130_fd_sc_hd__o21ai_2 _27386_ (.A1(_06622_),
    .A2(_06624_),
    .B1(_03331_),
    .Y(_03341_));
 sky130_fd_sc_hd__a211oi_2 _27387_ (.A1(_03337_),
    .A2(_03329_),
    .B1(_03336_),
    .C1(_03340_),
    .Y(_03342_));
 sky130_fd_sc_hd__nand3_1 _27388_ (.A(_03341_),
    .B(_03335_),
    .C(_03339_),
    .Y(_03343_));
 sky130_fd_sc_hd__o22a_1 _27389_ (.A1(_03067_),
    .A2(_03333_),
    .B1(_03338_),
    .B2(_03340_),
    .X(_03344_));
 sky130_fd_sc_hd__o22ai_2 _27390_ (.A1(_03067_),
    .A2(_03333_),
    .B1(_03338_),
    .B2(_03340_),
    .Y(_03346_));
 sky130_fd_sc_hd__o22ai_4 _27391_ (.A1(net141),
    .A2(net140),
    .B1(_03342_),
    .B2(_03344_),
    .Y(_03347_));
 sky130_fd_sc_hd__or3_1 _27392_ (.A(net141),
    .B(net140),
    .C(_03330_),
    .X(_03348_));
 sky130_fd_sc_hd__o211ai_4 _27393_ (.A1(net141),
    .A2(net140),
    .B1(_03343_),
    .C1(_03346_),
    .Y(_03349_));
 sky130_fd_sc_hd__o21ai_4 _27394_ (.A1(net131),
    .A2(_03330_),
    .B1(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__a211o_1 _27395_ (.A1(_03348_),
    .A2(_03349_),
    .B1(net137),
    .C1(net135),
    .X(_03351_));
 sky130_fd_sc_hd__a2bb2oi_2 _27396_ (.A1_N(net284),
    .A2_N(net281),
    .B1(_03348_),
    .B2(_03349_),
    .Y(_03352_));
 sky130_fd_sc_hd__o221ai_4 _27397_ (.A1(net284),
    .A2(net281),
    .B1(net131),
    .B2(_03331_),
    .C1(_03347_),
    .Y(_03353_));
 sky130_fd_sc_hd__o211a_1 _27398_ (.A1(net131),
    .A2(_03330_),
    .B1(_06314_),
    .C1(_03349_),
    .X(_03354_));
 sky130_fd_sc_hd__o2111ai_4 _27399_ (.A1(_03330_),
    .A2(net131),
    .B1(_06308_),
    .C1(_06306_),
    .D1(_03349_),
    .Y(_03355_));
 sky130_fd_sc_hd__a31oi_4 _27400_ (.A1(_02820_),
    .A2(_02837_),
    .A3(_03083_),
    .B1(_03081_),
    .Y(_03357_));
 sky130_fd_sc_hd__o21bai_2 _27401_ (.A1(_03352_),
    .A2(_03354_),
    .B1_N(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__nand3_1 _27402_ (.A(_03353_),
    .B(_03355_),
    .C(_03357_),
    .Y(_03359_));
 sky130_fd_sc_hd__a31oi_2 _27403_ (.A1(_03353_),
    .A2(_03357_),
    .A3(_03355_),
    .B1(_10953_),
    .Y(_03360_));
 sky130_fd_sc_hd__o211ai_1 _27404_ (.A1(net137),
    .A2(net135),
    .B1(_03358_),
    .C1(_03359_),
    .Y(_03361_));
 sky130_fd_sc_hd__a22oi_2 _27405_ (.A1(_10953_),
    .A2(_03350_),
    .B1(_03360_),
    .B2(_03358_),
    .Y(_03362_));
 sky130_fd_sc_hd__a32o_1 _27406_ (.A1(_10953_),
    .A2(_03332_),
    .A3(_03347_),
    .B1(_03360_),
    .B2(_03358_),
    .X(_03363_));
 sky130_fd_sc_hd__and3_1 _27407_ (.A(_11460_),
    .B(_11462_),
    .C(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__a2bb2oi_1 _27408_ (.A1_N(_06009_),
    .A2_N(net287),
    .B1(_03351_),
    .B2(_03361_),
    .Y(_03365_));
 sky130_fd_sc_hd__a21oi_1 _27409_ (.A1(_03360_),
    .A2(_03358_),
    .B1(_06014_),
    .Y(_03366_));
 sky130_fd_sc_hd__and3_1 _27410_ (.A(_03361_),
    .B(_06013_),
    .C(_03351_),
    .X(_03368_));
 sky130_fd_sc_hd__a221o_1 _27411_ (.A1(_10953_),
    .A2(_03350_),
    .B1(_03360_),
    .B2(_03358_),
    .C1(_06014_),
    .X(_03369_));
 sky130_fd_sc_hd__a21oi_1 _27412_ (.A1(_03351_),
    .A2(_03366_),
    .B1(_03365_),
    .Y(_03370_));
 sky130_fd_sc_hd__o22ai_1 _27413_ (.A1(_05767_),
    .A2(_03089_),
    .B1(_03106_),
    .B2(_03099_),
    .Y(_03371_));
 sky130_fd_sc_hd__o221ai_2 _27414_ (.A1(_05767_),
    .A2(_03089_),
    .B1(_03365_),
    .B2(_03368_),
    .C1(_03107_),
    .Y(_03372_));
 sky130_fd_sc_hd__nand3b_1 _27415_ (.A_N(_03365_),
    .B(_03371_),
    .C(_03369_),
    .Y(_03373_));
 sky130_fd_sc_hd__a31oi_1 _27416_ (.A1(_11465_),
    .A2(_03372_),
    .A3(_03373_),
    .B1(_03364_),
    .Y(_03374_));
 sky130_fd_sc_hd__nand3b_1 _27417_ (.A_N(_02553_),
    .B(_02556_),
    .C(_02254_),
    .Y(_03375_));
 sky130_fd_sc_hd__nor3_1 _27418_ (.A(_03375_),
    .B(_02852_),
    .C(_02851_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand2_1 _27419_ (.A(_03376_),
    .B(_03110_),
    .Y(_03377_));
 sky130_fd_sc_hd__o211ai_2 _27420_ (.A1(_03112_),
    .A2(_03109_),
    .B1(_03111_),
    .C1(_03377_),
    .Y(_03379_));
 sky130_fd_sc_hd__nand4_1 _27421_ (.A(_03376_),
    .B(_03111_),
    .C(_03110_),
    .D(_02256_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand2_1 _27422_ (.A(_03379_),
    .B(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__a311o_1 _27423_ (.A1(_11465_),
    .A2(_03372_),
    .A3(_03373_),
    .B1(_03364_),
    .C1(_05768_),
    .X(_03382_));
 sky130_fd_sc_hd__a21o_1 _27424_ (.A1(_05761_),
    .A2(_05764_),
    .B1(_03374_),
    .X(_03383_));
 sky130_fd_sc_hd__nand2_1 _27425_ (.A(_03382_),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__a21o_1 _27426_ (.A1(_03381_),
    .A2(_03384_),
    .B1(_11944_),
    .X(_03385_));
 sky130_fd_sc_hd__nand2_1 _27427_ (.A(_03385_),
    .B(_03374_),
    .Y(_03386_));
 sky130_fd_sc_hd__xnor2_1 _27428_ (.A(_03118_),
    .B(_03386_),
    .Y(net106));
 sky130_fd_sc_hd__or4_2 _27429_ (.A(_02562_),
    .B(_02856_),
    .C(_03115_),
    .D(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__a31o_1 _27430_ (.A1(_11471_),
    .A2(_03130_),
    .A3(_03135_),
    .B1(_06294_),
    .X(_03389_));
 sky130_fd_sc_hd__a311o_2 _27431_ (.A1(_11471_),
    .A2(_03130_),
    .A3(_03135_),
    .B1(net209),
    .C1(_06294_),
    .X(_03390_));
 sky130_fd_sc_hd__inv_2 _27432_ (.A(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__xor2_1 _27433_ (.A(_10970_),
    .B(_03389_),
    .X(_03392_));
 sky130_fd_sc_hd__xor2_1 _27434_ (.A(_10971_),
    .B(_03389_),
    .X(_03393_));
 sky130_fd_sc_hd__o21ai_2 _27435_ (.A1(_03141_),
    .A2(_03150_),
    .B1(_03392_),
    .Y(_03394_));
 sky130_fd_sc_hd__o211ai_2 _27436_ (.A1(net150),
    .A2(_03140_),
    .B1(_03151_),
    .C1(_03393_),
    .Y(_03395_));
 sky130_fd_sc_hd__nand3_2 _27437_ (.A(_03394_),
    .B(_03395_),
    .C(net209),
    .Y(_03396_));
 sky130_fd_sc_hd__o21a_1 _27438_ (.A1(net209),
    .A2(_03389_),
    .B1(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__and3_1 _27439_ (.A(_06904_),
    .B(_03390_),
    .C(_03396_),
    .X(_03398_));
 sky130_fd_sc_hd__a2bb2oi_1 _27440_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_03390_),
    .B2(_03396_),
    .Y(_03401_));
 sky130_fd_sc_hd__a2bb2o_2 _27441_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_03390_),
    .B2(_03396_),
    .X(_03402_));
 sky130_fd_sc_hd__a31o_1 _27442_ (.A1(_03394_),
    .A2(_03395_),
    .A3(net209),
    .B1(_10492_),
    .X(_03403_));
 sky130_fd_sc_hd__and3_1 _27443_ (.A(_03396_),
    .B(net150),
    .C(_03390_),
    .X(_03404_));
 sky130_fd_sc_hd__o2bb2ai_1 _27444_ (.A1_N(_03164_),
    .A2_N(_03166_),
    .B1(net152),
    .B2(_03155_),
    .Y(_03405_));
 sky130_fd_sc_hd__a31oi_2 _27445_ (.A1(_03164_),
    .A2(_03166_),
    .A3(_03172_),
    .B1(_03168_),
    .Y(_03406_));
 sky130_fd_sc_hd__o2111ai_4 _27446_ (.A1(_03403_),
    .A2(_03391_),
    .B1(_03172_),
    .C1(_03402_),
    .D1(_03405_),
    .Y(_03407_));
 sky130_fd_sc_hd__o21ai_2 _27447_ (.A1(_03401_),
    .A2(_03404_),
    .B1(_03406_),
    .Y(_03408_));
 sky130_fd_sc_hd__a21oi_1 _27448_ (.A1(_03407_),
    .A2(_03408_),
    .B1(_06904_),
    .Y(_03409_));
 sky130_fd_sc_hd__a21oi_1 _27449_ (.A1(_03390_),
    .A2(_03396_),
    .B1(_06903_),
    .Y(_03410_));
 sky130_fd_sc_hd__inv_2 _27450_ (.A(_03410_),
    .Y(_03412_));
 sky130_fd_sc_hd__nand3_2 _27451_ (.A(_03407_),
    .B(_03408_),
    .C(_06903_),
    .Y(_03413_));
 sky130_fd_sc_hd__a31o_1 _27452_ (.A1(_03407_),
    .A2(_03408_),
    .A3(_06903_),
    .B1(_03410_),
    .X(_03414_));
 sky130_fd_sc_hd__o31a_1 _27453_ (.A1(net229),
    .A2(net228),
    .A3(_03397_),
    .B1(_03413_),
    .X(_03415_));
 sky130_fd_sc_hd__a311o_2 _27454_ (.A1(_06904_),
    .A2(_03390_),
    .A3(_03396_),
    .B1(_07233_),
    .C1(_03409_),
    .X(_03416_));
 sky130_fd_sc_hd__inv_2 _27455_ (.A(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__and4_1 _27456_ (.A(_02368_),
    .B(_02369_),
    .C(_02664_),
    .D(_02666_),
    .X(_03418_));
 sky130_fd_sc_hd__nand3_1 _27457_ (.A(_03186_),
    .B(_03418_),
    .C(_02940_),
    .Y(_03419_));
 sky130_fd_sc_hd__o211ai_4 _27458_ (.A1(_03191_),
    .A2(_03185_),
    .B1(_03188_),
    .C1(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__nand4_1 _27459_ (.A(_03418_),
    .B(_02939_),
    .C(_02936_),
    .D(_02375_),
    .Y(_03421_));
 sky130_fd_sc_hd__nand3b_4 _27460_ (.A_N(_03421_),
    .B(_03188_),
    .C(_03186_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21oi_2 _27461_ (.A1(_03412_),
    .A2(_03413_),
    .B1(net152),
    .Y(_03424_));
 sky130_fd_sc_hd__a2bb2o_1 _27462_ (.A1_N(net170),
    .A2_N(net168),
    .B1(_03412_),
    .B2(_03413_),
    .X(_03425_));
 sky130_fd_sc_hd__o221a_1 _27463_ (.A1(net167),
    .A2(_10024_),
    .B1(_03397_),
    .B2(_06903_),
    .C1(_03413_),
    .X(_03426_));
 sky130_fd_sc_hd__a311o_2 _27464_ (.A1(_03407_),
    .A2(_03408_),
    .A3(_06903_),
    .B1(_03410_),
    .C1(net151),
    .X(_03427_));
 sky130_fd_sc_hd__nand4_2 _27465_ (.A(_03420_),
    .B(_03423_),
    .C(_03425_),
    .D(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__o2bb2ai_2 _27466_ (.A1_N(_03420_),
    .A2_N(_03423_),
    .B1(_03424_),
    .B2(_03426_),
    .Y(_03429_));
 sky130_fd_sc_hd__o211a_1 _27467_ (.A1(net207),
    .A2(net204),
    .B1(_03428_),
    .C1(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__o211ai_4 _27468_ (.A1(net207),
    .A2(net204),
    .B1(_03428_),
    .C1(_03429_),
    .Y(_03431_));
 sky130_fd_sc_hd__o211a_2 _27469_ (.A1(_03417_),
    .A2(_03430_),
    .B1(_07545_),
    .C1(_07547_),
    .X(_03432_));
 sky130_fd_sc_hd__a211o_1 _27470_ (.A1(_03416_),
    .A2(_03431_),
    .B1(_07544_),
    .C1(_07546_),
    .X(_03434_));
 sky130_fd_sc_hd__o311a_2 _27471_ (.A1(_07233_),
    .A2(_03398_),
    .A3(_03409_),
    .B1(_09594_),
    .C1(_03431_),
    .X(_03435_));
 sky130_fd_sc_hd__nand3_2 _27472_ (.A(_03431_),
    .B(_09594_),
    .C(_03416_),
    .Y(_03436_));
 sky130_fd_sc_hd__a21oi_1 _27473_ (.A1(_03416_),
    .A2(_03431_),
    .B1(_09594_),
    .Y(_03437_));
 sky130_fd_sc_hd__o22ai_4 _27474_ (.A1(net189),
    .A2(net186),
    .B1(_03417_),
    .B2(_03430_),
    .Y(_03438_));
 sky130_fd_sc_hd__a31o_1 _27475_ (.A1(_02954_),
    .A2(_03200_),
    .A3(_03206_),
    .B1(_03207_),
    .X(_03439_));
 sky130_fd_sc_hd__o22ai_2 _27476_ (.A1(_03183_),
    .A2(_03204_),
    .B1(_03207_),
    .B2(_03203_),
    .Y(_03440_));
 sky130_fd_sc_hd__o21bai_4 _27477_ (.A1(_03435_),
    .A2(_03437_),
    .B1_N(_03439_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand3_2 _27478_ (.A(_03436_),
    .B(_03438_),
    .C(_03439_),
    .Y(_03442_));
 sky130_fd_sc_hd__nand3_1 _27479_ (.A(_03441_),
    .B(_03442_),
    .C(_07548_),
    .Y(_03443_));
 sky130_fd_sc_hd__a31oi_2 _27480_ (.A1(_03441_),
    .A2(_03442_),
    .A3(_07548_),
    .B1(_03432_),
    .Y(_03445_));
 sky130_fd_sc_hd__a31o_1 _27481_ (.A1(_03441_),
    .A2(_03442_),
    .A3(_07548_),
    .B1(_03432_),
    .X(_03446_));
 sky130_fd_sc_hd__o311a_1 _27482_ (.A1(_08311_),
    .A2(net215),
    .A3(_02965_),
    .B1(_03220_),
    .C1(_03226_),
    .X(_03447_));
 sky130_fd_sc_hd__a22o_1 _27483_ (.A1(net178),
    .A2(_03219_),
    .B1(_03226_),
    .B2(_02967_),
    .X(_03448_));
 sky130_fd_sc_hd__o21ai_2 _27484_ (.A1(_03221_),
    .A2(_03227_),
    .B1(_03220_),
    .Y(_03449_));
 sky130_fd_sc_hd__a31oi_1 _27485_ (.A1(_03441_),
    .A2(_03442_),
    .A3(_07548_),
    .B1(_09140_),
    .Y(_03450_));
 sky130_fd_sc_hd__a31o_1 _27486_ (.A1(_03441_),
    .A2(_03442_),
    .A3(_07548_),
    .B1(_09140_),
    .X(_03451_));
 sky130_fd_sc_hd__a311oi_2 _27487_ (.A1(_03441_),
    .A2(_03442_),
    .A3(_07548_),
    .B1(_09140_),
    .C1(_03432_),
    .Y(_03452_));
 sky130_fd_sc_hd__a2bb2oi_4 _27488_ (.A1_N(net194),
    .A2_N(net191),
    .B1(_03434_),
    .B2(_03443_),
    .Y(_03453_));
 sky130_fd_sc_hd__o21ai_1 _27489_ (.A1(net194),
    .A2(net191),
    .B1(_03446_),
    .Y(_03454_));
 sky130_fd_sc_hd__a21oi_1 _27490_ (.A1(_03434_),
    .A2(_03450_),
    .B1(_03453_),
    .Y(_03456_));
 sky130_fd_sc_hd__o221ai_1 _27491_ (.A1(_03221_),
    .A2(_03447_),
    .B1(_03451_),
    .B2(_03432_),
    .C1(_03454_),
    .Y(_03457_));
 sky130_fd_sc_hd__o2bb2ai_1 _27492_ (.A1_N(_03220_),
    .A2_N(_03448_),
    .B1(_03452_),
    .B2(_03453_),
    .Y(_03458_));
 sky130_fd_sc_hd__nand3_1 _27493_ (.A(_03457_),
    .B(_03458_),
    .C(_07916_),
    .Y(_03459_));
 sky130_fd_sc_hd__a21oi_1 _27494_ (.A1(_03434_),
    .A2(_03443_),
    .B1(_07916_),
    .Y(_03460_));
 sky130_fd_sc_hd__inv_2 _27495_ (.A(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__o211ai_1 _27496_ (.A1(_03432_),
    .A2(_03451_),
    .B1(_03449_),
    .C1(_03454_),
    .Y(_03462_));
 sky130_fd_sc_hd__o22ai_1 _27497_ (.A1(_03221_),
    .A2(_03447_),
    .B1(_03452_),
    .B2(_03453_),
    .Y(_03463_));
 sky130_fd_sc_hd__nand3_2 _27498_ (.A(_03462_),
    .B(_03463_),
    .C(_07916_),
    .Y(_03464_));
 sky130_fd_sc_hd__o31a_2 _27499_ (.A1(net183),
    .A2(net182),
    .A3(_03445_),
    .B1(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__inv_2 _27500_ (.A(_03465_),
    .Y(_03467_));
 sky130_fd_sc_hd__o221a_2 _27501_ (.A1(_08293_),
    .A2(_08295_),
    .B1(_03445_),
    .B2(_07916_),
    .C1(_03464_),
    .X(_03468_));
 sky130_fd_sc_hd__o211ai_4 _27502_ (.A1(_03446_),
    .A2(_07916_),
    .B1(_08731_),
    .C1(_03459_),
    .Y(_03469_));
 sky130_fd_sc_hd__and3_1 _27503_ (.A(_03464_),
    .B(net178),
    .C(_03461_),
    .X(_03470_));
 sky130_fd_sc_hd__nand3_4 _27504_ (.A(_03464_),
    .B(net178),
    .C(_03461_),
    .Y(_03471_));
 sky130_fd_sc_hd__nand2_1 _27505_ (.A(_03469_),
    .B(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__o2bb2ai_1 _27506_ (.A1_N(_03121_),
    .A2_N(_03124_),
    .B1(_03236_),
    .B2(net201),
    .Y(_03473_));
 sky130_fd_sc_hd__nand3_4 _27507_ (.A(_03121_),
    .B(_03124_),
    .C(_03240_),
    .Y(_03474_));
 sky130_fd_sc_hd__a31oi_2 _27508_ (.A1(_03121_),
    .A2(_03124_),
    .A3(_03240_),
    .B1(_03237_),
    .Y(_03475_));
 sky130_fd_sc_hd__o2111ai_4 _27509_ (.A1(_03236_),
    .A2(net201),
    .B1(_03471_),
    .C1(_03469_),
    .D1(_03474_),
    .Y(_03476_));
 sky130_fd_sc_hd__a22o_2 _27510_ (.A1(_03469_),
    .A2(_03471_),
    .B1(_03474_),
    .B2(_03238_),
    .X(_03478_));
 sky130_fd_sc_hd__nand3_2 _27511_ (.A(_03478_),
    .B(net159),
    .C(_03476_),
    .Y(_03479_));
 sky130_fd_sc_hd__a22oi_2 _27512_ (.A1(_03469_),
    .A2(_03471_),
    .B1(_03473_),
    .B2(_03240_),
    .Y(_03480_));
 sky130_fd_sc_hd__o22ai_2 _27513_ (.A1(net181),
    .A2(net179),
    .B1(_03472_),
    .B2(_03475_),
    .Y(_03481_));
 sky130_fd_sc_hd__a31oi_4 _27514_ (.A1(_03478_),
    .A2(net159),
    .A3(_03476_),
    .B1(_03468_),
    .Y(_03482_));
 sky130_fd_sc_hd__a31o_1 _27515_ (.A1(_03478_),
    .A2(net159),
    .A3(_03476_),
    .B1(_03468_),
    .X(_03483_));
 sky130_fd_sc_hd__o211a_1 _27516_ (.A1(net159),
    .A2(_03467_),
    .B1(_03479_),
    .C1(net197),
    .X(_03484_));
 sky130_fd_sc_hd__o211ai_4 _27517_ (.A1(net159),
    .A2(_03467_),
    .B1(_03479_),
    .C1(net197),
    .Y(_03485_));
 sky130_fd_sc_hd__o221ai_4 _27518_ (.A1(net159),
    .A2(_03465_),
    .B1(_03480_),
    .B2(_03481_),
    .C1(net201),
    .Y(_03486_));
 sky130_fd_sc_hd__nand2_1 _27519_ (.A(_03485_),
    .B(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__o2111ai_2 _27520_ (.A1(_02439_),
    .A2(_02431_),
    .B1(_02437_),
    .C1(_02735_),
    .D1(_02736_),
    .Y(_03489_));
 sky130_fd_sc_hd__a21oi_1 _27521_ (.A1(_07565_),
    .A2(_02991_),
    .B1(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__nor3_1 _27522_ (.A(_02996_),
    .B(_03489_),
    .C(_02998_),
    .Y(_03491_));
 sky130_fd_sc_hd__o211ai_2 _27523_ (.A1(_07565_),
    .A2(_02991_),
    .B1(_03490_),
    .C1(_03255_),
    .Y(_03492_));
 sky130_fd_sc_hd__o211ai_4 _27524_ (.A1(_03261_),
    .A2(_03254_),
    .B1(_03257_),
    .C1(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__nand4_4 _27525_ (.A(_03491_),
    .B(_03257_),
    .C(_03255_),
    .D(_02451_),
    .Y(_03494_));
 sky130_fd_sc_hd__nand2_1 _27526_ (.A(_03493_),
    .B(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__a21oi_2 _27527_ (.A1(_03493_),
    .A2(_03494_),
    .B1(_03487_),
    .Y(_03496_));
 sky130_fd_sc_hd__a31o_1 _27528_ (.A1(_03487_),
    .A2(_03493_),
    .A3(_03494_),
    .B1(_08715_),
    .X(_03497_));
 sky130_fd_sc_hd__and3_1 _27529_ (.A(_03482_),
    .B(_08713_),
    .C(_08710_),
    .X(_03498_));
 sky130_fd_sc_hd__a311o_1 _27530_ (.A1(_03478_),
    .A2(net159),
    .A3(_03476_),
    .B1(net149),
    .C1(_03468_),
    .X(_03500_));
 sky130_fd_sc_hd__a22o_1 _27531_ (.A1(_03485_),
    .A2(_03486_),
    .B1(_03493_),
    .B2(_03494_),
    .X(_03501_));
 sky130_fd_sc_hd__o211ai_4 _27532_ (.A1(_03482_),
    .A2(net197),
    .B1(_03494_),
    .C1(_03493_),
    .Y(_03502_));
 sky130_fd_sc_hd__o2111ai_4 _27533_ (.A1(net197),
    .A2(_03482_),
    .B1(_03485_),
    .C1(_03493_),
    .D1(_03494_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand3_2 _27534_ (.A(_03501_),
    .B(_03503_),
    .C(net149),
    .Y(_03504_));
 sky130_fd_sc_hd__a31o_1 _27535_ (.A1(_03501_),
    .A2(_03503_),
    .A3(net149),
    .B1(_03498_),
    .X(_03505_));
 sky130_fd_sc_hd__o221a_1 _27536_ (.A1(net149),
    .A2(_03482_),
    .B1(_03496_),
    .B2(_03497_),
    .C1(_09124_),
    .X(_03506_));
 sky130_fd_sc_hd__a211o_2 _27537_ (.A1(_03500_),
    .A2(_03504_),
    .B1(net148),
    .C1(net147),
    .X(_03507_));
 sky130_fd_sc_hd__a311oi_4 _27538_ (.A1(_03501_),
    .A2(_03503_),
    .A3(net149),
    .B1(_03498_),
    .C1(_07936_),
    .Y(_03508_));
 sky130_fd_sc_hd__nand3_4 _27539_ (.A(_03504_),
    .B(_07935_),
    .C(_03500_),
    .Y(_03509_));
 sky130_fd_sc_hd__o221ai_4 _27540_ (.A1(net149),
    .A2(_03482_),
    .B1(_03496_),
    .B2(_03497_),
    .C1(_07936_),
    .Y(_03512_));
 sky130_fd_sc_hd__o211a_1 _27541_ (.A1(_07246_),
    .A2(_03010_),
    .B1(_03022_),
    .C1(_03280_),
    .X(_03513_));
 sky130_fd_sc_hd__o211a_1 _27542_ (.A1(_03009_),
    .A2(net223),
    .B1(_03277_),
    .C1(_03273_),
    .X(_03514_));
 sky130_fd_sc_hd__a31o_1 _27543_ (.A1(_03013_),
    .A2(_03273_),
    .A3(_03277_),
    .B1(_03279_),
    .X(_03515_));
 sky130_fd_sc_hd__a21oi_1 _27544_ (.A1(_03274_),
    .A2(_03277_),
    .B1(_03279_),
    .Y(_03516_));
 sky130_fd_sc_hd__a21oi_2 _27545_ (.A1(_03509_),
    .A2(_03512_),
    .B1(_03515_),
    .Y(_03517_));
 sky130_fd_sc_hd__o2bb2ai_1 _27546_ (.A1_N(_03509_),
    .A2_N(_03512_),
    .B1(_03513_),
    .B2(_03276_),
    .Y(_03518_));
 sky130_fd_sc_hd__o211a_1 _27547_ (.A1(_03279_),
    .A2(_03514_),
    .B1(_03512_),
    .C1(_03509_),
    .X(_03519_));
 sky130_fd_sc_hd__nand3_1 _27548_ (.A(_03509_),
    .B(_03515_),
    .C(_03512_),
    .Y(_03520_));
 sky130_fd_sc_hd__a31oi_1 _27549_ (.A1(_03509_),
    .A2(_03515_),
    .A3(_03512_),
    .B1(_09124_),
    .Y(_03521_));
 sky130_fd_sc_hd__o21ai_2 _27550_ (.A1(net148),
    .A2(net147),
    .B1(_03520_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand3_1 _27551_ (.A(net145),
    .B(_03518_),
    .C(_03520_),
    .Y(_03524_));
 sky130_fd_sc_hd__o22ai_2 _27552_ (.A1(net148),
    .A2(net147),
    .B1(_03517_),
    .B2(_03519_),
    .Y(_03525_));
 sky130_fd_sc_hd__a221o_1 _27553_ (.A1(_09124_),
    .A2(_03505_),
    .B1(_03521_),
    .B2(_03518_),
    .C1(net144),
    .X(_03526_));
 sky130_fd_sc_hd__o211ai_4 _27554_ (.A1(_03026_),
    .A2(_06922_),
    .B1(_03294_),
    .C1(_03044_),
    .Y(_03527_));
 sky130_fd_sc_hd__a31oi_2 _27555_ (.A1(_03028_),
    .A2(_03044_),
    .A3(_03294_),
    .B1(_03291_),
    .Y(_03528_));
 sky130_fd_sc_hd__a31o_1 _27556_ (.A1(_03028_),
    .A2(_03044_),
    .A3(_03294_),
    .B1(_03291_),
    .X(_03529_));
 sky130_fd_sc_hd__o21ai_1 _27557_ (.A1(_03517_),
    .A2(_03523_),
    .B1(_07564_),
    .Y(_03530_));
 sky130_fd_sc_hd__a211oi_1 _27558_ (.A1(_03521_),
    .A2(_03518_),
    .B1(_03506_),
    .C1(_07565_),
    .Y(_03531_));
 sky130_fd_sc_hd__o211ai_4 _27559_ (.A1(_03517_),
    .A2(_03523_),
    .B1(_07564_),
    .C1(_03507_),
    .Y(_03532_));
 sky130_fd_sc_hd__a2bb2oi_2 _27560_ (.A1_N(net221),
    .A2_N(net219),
    .B1(_03507_),
    .B2(_03524_),
    .Y(_03534_));
 sky130_fd_sc_hd__o221ai_4 _27561_ (.A1(net221),
    .A2(net219),
    .B1(net145),
    .B2(_03505_),
    .C1(_03525_),
    .Y(_03535_));
 sky130_fd_sc_hd__o211ai_1 _27562_ (.A1(_03506_),
    .A2(_03530_),
    .B1(_03535_),
    .C1(_03529_),
    .Y(_03536_));
 sky130_fd_sc_hd__o21ai_1 _27563_ (.A1(_03531_),
    .A2(_03534_),
    .B1(_03528_),
    .Y(_03537_));
 sky130_fd_sc_hd__o211ai_2 _27564_ (.A1(net156),
    .A2(net154),
    .B1(_03536_),
    .C1(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__a211o_2 _27565_ (.A1(_03507_),
    .A2(_03524_),
    .B1(net156),
    .C1(net154),
    .X(_03539_));
 sky130_fd_sc_hd__o2111ai_4 _27566_ (.A1(net223),
    .A2(_03288_),
    .B1(_03527_),
    .C1(_03532_),
    .D1(_03535_),
    .Y(_03540_));
 sky130_fd_sc_hd__o2bb2ai_1 _27567_ (.A1_N(_03292_),
    .A2_N(_03527_),
    .B1(_03531_),
    .B2(_03534_),
    .Y(_03541_));
 sky130_fd_sc_hd__o211ai_4 _27568_ (.A1(net156),
    .A2(net154),
    .B1(_03540_),
    .C1(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__nand2_1 _27569_ (.A(_03539_),
    .B(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__o211ai_4 _27570_ (.A1(_07242_),
    .A2(net248),
    .B1(_03526_),
    .C1(_03538_),
    .Y(_03545_));
 sky130_fd_sc_hd__and3_1 _27571_ (.A(_03542_),
    .B(_07246_),
    .C(_03539_),
    .X(_03546_));
 sky130_fd_sc_hd__o211ai_4 _27572_ (.A1(_07244_),
    .A2(net247),
    .B1(_03539_),
    .C1(_03542_),
    .Y(_03547_));
 sky130_fd_sc_hd__nand2_2 _27573_ (.A(_03545_),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__o22ai_1 _27574_ (.A1(_06922_),
    .A2(_03305_),
    .B1(_03325_),
    .B2(_03316_),
    .Y(_03549_));
 sky130_fd_sc_hd__a2bb2oi_2 _27575_ (.A1_N(_06922_),
    .A2_N(_03305_),
    .B1(_03317_),
    .B2(_03324_),
    .Y(_03550_));
 sky130_fd_sc_hd__a21oi_1 _27576_ (.A1(_03549_),
    .A2(_03548_),
    .B1(_09578_),
    .Y(_03551_));
 sky130_fd_sc_hd__o21ai_1 _27577_ (.A1(_03548_),
    .A2(_03549_),
    .B1(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__a22o_2 _27578_ (.A1(_09575_),
    .A2(_09577_),
    .B1(_03539_),
    .B2(_03542_),
    .X(_03553_));
 sky130_fd_sc_hd__o311a_2 _27579_ (.A1(_06918_),
    .A2(net249),
    .A3(_03305_),
    .B1(_03326_),
    .C1(_03548_),
    .X(_03554_));
 sky130_fd_sc_hd__o21ai_4 _27580_ (.A1(_03548_),
    .A2(_03550_),
    .B1(net132),
    .Y(_03556_));
 sky130_fd_sc_hd__a31o_1 _27581_ (.A1(_03307_),
    .A2(_03326_),
    .A3(_03548_),
    .B1(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__o21ai_4 _27582_ (.A1(_03554_),
    .A2(_03556_),
    .B1(_03553_),
    .Y(_03558_));
 sky130_fd_sc_hd__o2bb2a_2 _27583_ (.A1_N(_09578_),
    .A2_N(_03543_),
    .B1(_03554_),
    .B2(_03556_),
    .X(_03559_));
 sky130_fd_sc_hd__o211ai_4 _27584_ (.A1(_03543_),
    .A2(net132),
    .B1(net226),
    .C1(_03552_),
    .Y(_03560_));
 sky130_fd_sc_hd__inv_2 _27585_ (.A(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__and3_1 _27586_ (.A(_03557_),
    .B(_06922_),
    .C(_03553_),
    .X(_03562_));
 sky130_fd_sc_hd__o211ai_4 _27587_ (.A1(_03554_),
    .A2(_03556_),
    .B1(_06922_),
    .C1(_03553_),
    .Y(_03563_));
 sky130_fd_sc_hd__nand2_1 _27588_ (.A(_03560_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__and4_1 _27589_ (.A(_02512_),
    .B(_02514_),
    .C(_02807_),
    .D(_02809_),
    .X(_03565_));
 sky130_fd_sc_hd__o211a_1 _27590_ (.A1(_03049_),
    .A2(_03066_),
    .B1(_03565_),
    .C1(_03071_),
    .X(_03567_));
 sky130_fd_sc_hd__o211ai_1 _27591_ (.A1(_03049_),
    .A2(_03066_),
    .B1(_03565_),
    .C1(_03071_),
    .Y(_03568_));
 sky130_fd_sc_hd__a31oi_2 _27592_ (.A1(_03328_),
    .A2(_03329_),
    .A3(_06629_),
    .B1(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _27593_ (.A(_03339_),
    .B(_03567_),
    .Y(_03570_));
 sky130_fd_sc_hd__o211a_1 _27594_ (.A1(_03336_),
    .A2(_03338_),
    .B1(_03341_),
    .C1(_03570_),
    .X(_03571_));
 sky130_fd_sc_hd__o211ai_4 _27595_ (.A1(_03336_),
    .A2(_03338_),
    .B1(_03341_),
    .C1(_03570_),
    .Y(_03572_));
 sky130_fd_sc_hd__nand4_1 _27596_ (.A(_02523_),
    .B(_03068_),
    .C(_03071_),
    .D(_03565_),
    .Y(_03573_));
 sky130_fd_sc_hd__o211ai_4 _27597_ (.A1(_06629_),
    .A2(_03330_),
    .B1(_02523_),
    .C1(_03569_),
    .Y(_03574_));
 sky130_fd_sc_hd__a31o_2 _27598_ (.A1(_02523_),
    .A2(_03341_),
    .A3(_03569_),
    .B1(_03571_),
    .X(_03575_));
 sky130_fd_sc_hd__a21oi_1 _27599_ (.A1(_03572_),
    .A2(_03574_),
    .B1(_03564_),
    .Y(_03576_));
 sky130_fd_sc_hd__a21o_1 _27600_ (.A1(_03572_),
    .A2(_03574_),
    .B1(_03564_),
    .X(_03578_));
 sky130_fd_sc_hd__a31oi_1 _27601_ (.A1(_03564_),
    .A2(_03572_),
    .A3(_03574_),
    .B1(_10479_),
    .Y(_03579_));
 sky130_fd_sc_hd__a31o_1 _27602_ (.A1(_03564_),
    .A2(_03572_),
    .A3(_03574_),
    .B1(_10479_),
    .X(_03580_));
 sky130_fd_sc_hd__or3_1 _27603_ (.A(net141),
    .B(net140),
    .C(_03559_),
    .X(_03581_));
 sky130_fd_sc_hd__a22oi_1 _27604_ (.A1(_03560_),
    .A2(_03563_),
    .B1(_03572_),
    .B2(_03574_),
    .Y(_03582_));
 sky130_fd_sc_hd__a22o_1 _27605_ (.A1(_03560_),
    .A2(_03563_),
    .B1(_03572_),
    .B2(_03574_),
    .X(_03583_));
 sky130_fd_sc_hd__o31ai_1 _27606_ (.A1(_03573_),
    .A2(_03340_),
    .A3(_03338_),
    .B1(_03563_),
    .Y(_03584_));
 sky130_fd_sc_hd__o211ai_4 _27607_ (.A1(_03558_),
    .A2(net226),
    .B1(_03574_),
    .C1(_03572_),
    .Y(_03585_));
 sky130_fd_sc_hd__o2111a_1 _27608_ (.A1(net226),
    .A2(_03558_),
    .B1(_03560_),
    .C1(_03572_),
    .D1(_03574_),
    .X(_03586_));
 sky130_fd_sc_hd__o221ai_4 _27609_ (.A1(net141),
    .A2(net140),
    .B1(_03561_),
    .B2(_03585_),
    .C1(_03583_),
    .Y(_03587_));
 sky130_fd_sc_hd__a32o_2 _27610_ (.A1(_10479_),
    .A2(_03553_),
    .A3(_03557_),
    .B1(_03579_),
    .B2(_03578_),
    .X(_03589_));
 sky130_fd_sc_hd__inv_2 _27611_ (.A(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__o311a_2 _27612_ (.A1(_10479_),
    .A2(_03582_),
    .A3(_03586_),
    .B1(_03581_),
    .C1(_06629_),
    .X(_03591_));
 sky130_fd_sc_hd__nand3_4 _27613_ (.A(_03587_),
    .B(_06629_),
    .C(_03581_),
    .Y(_03592_));
 sky130_fd_sc_hd__a221oi_2 _27614_ (.A1(_10479_),
    .A2(_03559_),
    .B1(_03579_),
    .B2(_03578_),
    .C1(_06629_),
    .Y(_03593_));
 sky130_fd_sc_hd__o221ai_4 _27615_ (.A1(net131),
    .A2(_03558_),
    .B1(_03576_),
    .B2(_03580_),
    .C1(_06630_),
    .Y(_03594_));
 sky130_fd_sc_hd__a21oi_1 _27616_ (.A1(_06315_),
    .A2(_03350_),
    .B1(_03357_),
    .Y(_03595_));
 sky130_fd_sc_hd__a31o_1 _27617_ (.A1(_06315_),
    .A2(_03332_),
    .A3(_03347_),
    .B1(_03357_),
    .X(_03596_));
 sky130_fd_sc_hd__o32a_1 _27618_ (.A1(net284),
    .A2(net281),
    .A3(_03350_),
    .B1(_03352_),
    .B2(_03357_),
    .X(_03597_));
 sky130_fd_sc_hd__a21oi_2 _27619_ (.A1(_03357_),
    .A2(_03355_),
    .B1(_03352_),
    .Y(_03598_));
 sky130_fd_sc_hd__a21oi_1 _27620_ (.A1(_03592_),
    .A2(_03594_),
    .B1(_03597_),
    .Y(_03600_));
 sky130_fd_sc_hd__o2bb2ai_1 _27621_ (.A1_N(_03592_),
    .A2_N(_03594_),
    .B1(_03595_),
    .B2(_03354_),
    .Y(_03601_));
 sky130_fd_sc_hd__o2111a_1 _27622_ (.A1(_03350_),
    .A2(_06315_),
    .B1(_03594_),
    .C1(_03592_),
    .D1(_03596_),
    .X(_03602_));
 sky130_fd_sc_hd__o311ai_4 _27623_ (.A1(_03598_),
    .A2(_03593_),
    .A3(_03591_),
    .B1(_10954_),
    .C1(_03601_),
    .Y(_03603_));
 sky130_fd_sc_hd__o22ai_2 _27624_ (.A1(net137),
    .A2(net135),
    .B1(_03600_),
    .B2(_03602_),
    .Y(_03604_));
 sky130_fd_sc_hd__o31a_1 _27625_ (.A1(net137),
    .A2(net135),
    .A3(_03589_),
    .B1(_03603_),
    .X(_03605_));
 sky130_fd_sc_hd__o31a_1 _27626_ (.A1(net137),
    .A2(net135),
    .A3(_03590_),
    .B1(_03604_),
    .X(_03606_));
 sky130_fd_sc_hd__o221ai_4 _27627_ (.A1(_05767_),
    .A2(_03089_),
    .B1(_03362_),
    .B2(_06013_),
    .C1(_03107_),
    .Y(_03607_));
 sky130_fd_sc_hd__o211ai_4 _27628_ (.A1(_10954_),
    .A2(_03589_),
    .B1(_06314_),
    .C1(_03603_),
    .Y(_03608_));
 sky130_fd_sc_hd__o221ai_4 _27629_ (.A1(net284),
    .A2(net281),
    .B1(_10954_),
    .B2(_03590_),
    .C1(_03604_),
    .Y(_03609_));
 sky130_fd_sc_hd__o2111a_1 _27630_ (.A1(_06014_),
    .A2(_03363_),
    .B1(_03607_),
    .C1(_03608_),
    .D1(_03609_),
    .X(_03611_));
 sky130_fd_sc_hd__a22oi_1 _27631_ (.A1(_03369_),
    .A2(_03607_),
    .B1(_03608_),
    .B2(_03609_),
    .Y(_03612_));
 sky130_fd_sc_hd__o21ai_1 _27632_ (.A1(_03611_),
    .A2(_03612_),
    .B1(_11465_),
    .Y(_03613_));
 sky130_fd_sc_hd__or3_1 _27633_ (.A(_11459_),
    .B(net129),
    .C(_03605_),
    .X(_03614_));
 sky130_fd_sc_hd__o21a_1 _27634_ (.A1(_11465_),
    .A2(_03606_),
    .B1(_03613_),
    .X(_03615_));
 sky130_fd_sc_hd__o31a_1 _27635_ (.A1(_11464_),
    .A2(_03611_),
    .A3(_03612_),
    .B1(_06013_),
    .X(_03616_));
 sky130_fd_sc_hd__o21ai_1 _27636_ (.A1(_11465_),
    .A2(_03605_),
    .B1(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__o211ai_2 _27637_ (.A1(_11465_),
    .A2(_03606_),
    .B1(_03613_),
    .C1(_06014_),
    .Y(_03618_));
 sky130_fd_sc_hd__nand2_1 _27638_ (.A(_03617_),
    .B(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__nand3_1 _27639_ (.A(_03379_),
    .B(_03380_),
    .C(_03382_),
    .Y(_03620_));
 sky130_fd_sc_hd__a31oi_1 _27640_ (.A1(_03383_),
    .A2(_03619_),
    .A3(_03620_),
    .B1(_11944_),
    .Y(_03623_));
 sky130_fd_sc_hd__or2_1 _27641_ (.A(_03615_),
    .B(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__and3_1 _27642_ (.A(_05119_),
    .B(_03387_),
    .C(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__a21oi_1 _27643_ (.A1(_05119_),
    .A2(_03387_),
    .B1(_03624_),
    .Y(_03626_));
 sky130_fd_sc_hd__nor2_1 _27644_ (.A(_03625_),
    .B(_03626_),
    .Y(net107));
 sky130_fd_sc_hd__or4_1 _27645_ (.A(_02859_),
    .B(_03115_),
    .C(_03386_),
    .D(_03624_),
    .X(_03627_));
 sky130_fd_sc_hd__o32a_1 _27646_ (.A1(_03399_),
    .A2(net24),
    .A3(_10962_),
    .B1(_10970_),
    .B2(_03389_),
    .X(_03628_));
 sky130_fd_sc_hd__nand2_1 _27647_ (.A(_03394_),
    .B(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__a22o_1 _27648_ (.A1(_06609_),
    .A2(_06611_),
    .B1(_03394_),
    .B2(_03628_),
    .X(_03630_));
 sky130_fd_sc_hd__or3_4 _27649_ (.A(net229),
    .B(net228),
    .C(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__and3_1 _27650_ (.A(_03629_),
    .B(net209),
    .C(_10971_),
    .X(_03633_));
 sky130_fd_sc_hd__a211o_1 _27651_ (.A1(_03394_),
    .A2(_03628_),
    .B1(_06613_),
    .C1(_10970_),
    .X(_03634_));
 sky130_fd_sc_hd__a22o_1 _27652_ (.A1(_10966_),
    .A2(_10968_),
    .B1(_03629_),
    .B2(net209),
    .X(_03635_));
 sky130_fd_sc_hd__and2_1 _27653_ (.A(_03634_),
    .B(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__nand2_1 _27654_ (.A(_03634_),
    .B(_03635_),
    .Y(_03637_));
 sky130_fd_sc_hd__o21ai_1 _27655_ (.A1(_03404_),
    .A2(_03406_),
    .B1(_03402_),
    .Y(_03638_));
 sky130_fd_sc_hd__a21oi_4 _27656_ (.A1(_03402_),
    .A2(_03407_),
    .B1(_03637_),
    .Y(_03639_));
 sky130_fd_sc_hd__nand2_1 _27657_ (.A(_03638_),
    .B(_03636_),
    .Y(_03640_));
 sky130_fd_sc_hd__o211ai_2 _27658_ (.A1(_03404_),
    .A2(_03406_),
    .B1(_03637_),
    .C1(_03402_),
    .Y(_03641_));
 sky130_fd_sc_hd__o21ai_4 _27659_ (.A1(net229),
    .A2(net228),
    .B1(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__o211ai_1 _27660_ (.A1(net229),
    .A2(net228),
    .B1(_03640_),
    .C1(_03641_),
    .Y(_03644_));
 sky130_fd_sc_hd__o21ai_4 _27661_ (.A1(_03642_),
    .A2(_03639_),
    .B1(_03631_),
    .Y(_03645_));
 sky130_fd_sc_hd__a211o_1 _27662_ (.A1(_03631_),
    .A2(_03644_),
    .B1(net207),
    .C1(net204),
    .X(_03646_));
 sky130_fd_sc_hd__o21ai_2 _27663_ (.A1(_10487_),
    .A2(net165),
    .B1(_03645_),
    .Y(_03647_));
 sky130_fd_sc_hd__and3_1 _27664_ (.A(_03644_),
    .B(net150),
    .C(_03631_),
    .X(_03648_));
 sky130_fd_sc_hd__o211ai_4 _27665_ (.A1(_03642_),
    .A2(_03639_),
    .B1(_03631_),
    .C1(net150),
    .Y(_03649_));
 sky130_fd_sc_hd__nand2_1 _27666_ (.A(_03647_),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__o2bb2ai_2 _27667_ (.A1_N(_03420_),
    .A2_N(_03423_),
    .B1(net152),
    .B2(_03415_),
    .Y(_03651_));
 sky130_fd_sc_hd__a31oi_4 _27668_ (.A1(_03420_),
    .A2(_03423_),
    .A3(_03427_),
    .B1(_03424_),
    .Y(_03652_));
 sky130_fd_sc_hd__a22oi_4 _27669_ (.A1(_03647_),
    .A2(_03649_),
    .B1(_03651_),
    .B2(_03427_),
    .Y(_03653_));
 sky130_fd_sc_hd__nand2_1 _27670_ (.A(_03650_),
    .B(_03652_),
    .Y(_03655_));
 sky130_fd_sc_hd__o2111a_1 _27671_ (.A1(net151),
    .A2(_03414_),
    .B1(_03647_),
    .C1(_03649_),
    .D1(_03651_),
    .X(_03656_));
 sky130_fd_sc_hd__o211ai_2 _27672_ (.A1(_03650_),
    .A2(_03652_),
    .B1(_03655_),
    .C1(_07233_),
    .Y(_03657_));
 sky130_fd_sc_hd__o22ai_4 _27673_ (.A1(net207),
    .A2(net204),
    .B1(_03653_),
    .B2(_03656_),
    .Y(_03658_));
 sky130_fd_sc_hd__o31a_1 _27674_ (.A1(_07232_),
    .A2(_03653_),
    .A3(_03656_),
    .B1(_03646_),
    .X(_03659_));
 sky130_fd_sc_hd__o311a_2 _27675_ (.A1(net207),
    .A2(_03645_),
    .A3(net204),
    .B1(_07550_),
    .C1(_03658_),
    .X(_03660_));
 sky130_fd_sc_hd__or3_2 _27676_ (.A(_07544_),
    .B(_07546_),
    .C(_03659_),
    .X(_03661_));
 sky130_fd_sc_hd__o311a_1 _27677_ (.A1(net207),
    .A2(_03645_),
    .A3(net204),
    .B1(net151),
    .C1(_03658_),
    .X(_03662_));
 sky130_fd_sc_hd__o221ai_4 _27678_ (.A1(net170),
    .A2(net168),
    .B1(_03645_),
    .B2(_07233_),
    .C1(_03658_),
    .Y(_03663_));
 sky130_fd_sc_hd__o211ai_4 _27679_ (.A1(net167),
    .A2(_10024_),
    .B1(_03646_),
    .C1(_03657_),
    .Y(_03664_));
 sky130_fd_sc_hd__and4_1 _27680_ (.A(_02679_),
    .B(_02680_),
    .C(_02952_),
    .D(_02954_),
    .X(_03666_));
 sky130_fd_sc_hd__nand3_1 _27681_ (.A(_03209_),
    .B(_03436_),
    .C(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__o211ai_4 _27682_ (.A1(_03440_),
    .A2(_03435_),
    .B1(_03438_),
    .C1(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__and4_1 _27683_ (.A(_03666_),
    .B(_03208_),
    .C(_03206_),
    .D(_02688_),
    .X(_03669_));
 sky130_fd_sc_hd__nand3_4 _27684_ (.A(_03669_),
    .B(_03438_),
    .C(_03436_),
    .Y(_03670_));
 sky130_fd_sc_hd__a22o_2 _27685_ (.A1(_03663_),
    .A2(_03664_),
    .B1(_03668_),
    .B2(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__nand3_2 _27686_ (.A(_03664_),
    .B(_03668_),
    .C(_03670_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand4_4 _27687_ (.A(_03663_),
    .B(_03664_),
    .C(_03668_),
    .D(_03670_),
    .Y(_03673_));
 sky130_fd_sc_hd__o221a_1 _27688_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_03662_),
    .B2(_03672_),
    .C1(_03671_),
    .X(_03674_));
 sky130_fd_sc_hd__nand3_2 _27689_ (.A(_03671_),
    .B(_03673_),
    .C(_07548_),
    .Y(_03675_));
 sky130_fd_sc_hd__a2bb2o_2 _27690_ (.A1_N(_07909_),
    .A2_N(_07911_),
    .B1(_03661_),
    .B2(_03675_),
    .X(_03677_));
 sky130_fd_sc_hd__inv_2 _27691_ (.A(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__a31o_1 _27692_ (.A1(_03671_),
    .A2(_03673_),
    .A3(_07548_),
    .B1(net171),
    .X(_03679_));
 sky130_fd_sc_hd__a311oi_4 _27693_ (.A1(_03671_),
    .A2(_03673_),
    .A3(_07548_),
    .B1(net171),
    .C1(_03660_),
    .Y(_03680_));
 sky130_fd_sc_hd__nand3_2 _27694_ (.A(_03675_),
    .B(_09594_),
    .C(_03661_),
    .Y(_03681_));
 sky130_fd_sc_hd__a2bb2oi_2 _27695_ (.A1_N(net189),
    .A2_N(net186),
    .B1(_03661_),
    .B2(_03675_),
    .Y(_03682_));
 sky130_fd_sc_hd__o22ai_4 _27696_ (.A1(net189),
    .A2(net186),
    .B1(_03660_),
    .B2(_03674_),
    .Y(_03683_));
 sky130_fd_sc_hd__o32a_1 _27697_ (.A1(net194),
    .A2(net191),
    .A3(_03446_),
    .B1(_03449_),
    .B2(_03453_),
    .X(_03684_));
 sky130_fd_sc_hd__o22ai_4 _27698_ (.A1(_03432_),
    .A2(_03451_),
    .B1(_03453_),
    .B2(_03449_),
    .Y(_03685_));
 sky130_fd_sc_hd__o21ai_4 _27699_ (.A1(_03680_),
    .A2(_03682_),
    .B1(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__o211ai_4 _27700_ (.A1(_03660_),
    .A2(_03679_),
    .B1(_03684_),
    .C1(_03683_),
    .Y(_03688_));
 sky130_fd_sc_hd__o311a_1 _27701_ (.A1(_03680_),
    .A2(_03682_),
    .A3(_03685_),
    .B1(_07916_),
    .C1(_03686_),
    .X(_03689_));
 sky130_fd_sc_hd__nand3_2 _27702_ (.A(_03686_),
    .B(_03688_),
    .C(_07916_),
    .Y(_03690_));
 sky130_fd_sc_hd__a31o_2 _27703_ (.A1(_03686_),
    .A2(_03688_),
    .A3(_07916_),
    .B1(_03678_),
    .X(_03691_));
 sky130_fd_sc_hd__o311a_1 _27704_ (.A1(_08311_),
    .A2(net215),
    .A3(_03236_),
    .B1(_03469_),
    .C1(_03474_),
    .X(_03692_));
 sky130_fd_sc_hd__o21ai_1 _27705_ (.A1(net178),
    .A2(_03465_),
    .B1(_03475_),
    .Y(_03693_));
 sky130_fd_sc_hd__a22o_1 _27706_ (.A1(_03465_),
    .A2(net178),
    .B1(_03238_),
    .B2(_03474_),
    .X(_03694_));
 sky130_fd_sc_hd__a31oi_2 _27707_ (.A1(_03238_),
    .A2(_03469_),
    .A3(_03474_),
    .B1(_03470_),
    .Y(_03695_));
 sky130_fd_sc_hd__a31oi_1 _27708_ (.A1(_03686_),
    .A2(_03688_),
    .A3(_07916_),
    .B1(_09140_),
    .Y(_03696_));
 sky130_fd_sc_hd__a311oi_4 _27709_ (.A1(_03686_),
    .A2(_03688_),
    .A3(_07916_),
    .B1(_09140_),
    .C1(_03678_),
    .Y(_03697_));
 sky130_fd_sc_hd__nand3_2 _27710_ (.A(_03690_),
    .B(_09139_),
    .C(_03677_),
    .Y(_03699_));
 sky130_fd_sc_hd__a2bb2oi_2 _27711_ (.A1_N(net194),
    .A2_N(net191),
    .B1(_03677_),
    .B2(_03690_),
    .Y(_03700_));
 sky130_fd_sc_hd__o22ai_2 _27712_ (.A1(net194),
    .A2(net191),
    .B1(_03678_),
    .B2(_03689_),
    .Y(_03701_));
 sky130_fd_sc_hd__a21oi_1 _27713_ (.A1(_03677_),
    .A2(_03696_),
    .B1(_03700_),
    .Y(_03702_));
 sky130_fd_sc_hd__o211ai_2 _27714_ (.A1(_03470_),
    .A2(_03692_),
    .B1(_03699_),
    .C1(_03701_),
    .Y(_03703_));
 sky130_fd_sc_hd__o2bb2ai_1 _27715_ (.A1_N(_03469_),
    .A2_N(_03694_),
    .B1(_03697_),
    .B2(_03700_),
    .Y(_03704_));
 sky130_fd_sc_hd__o211ai_4 _27716_ (.A1(net181),
    .A2(net179),
    .B1(_03703_),
    .C1(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__a211o_1 _27717_ (.A1(_03677_),
    .A2(_03690_),
    .B1(net181),
    .C1(net179),
    .X(_03706_));
 sky130_fd_sc_hd__nand3_1 _27718_ (.A(_03701_),
    .B(_03695_),
    .C(_03699_),
    .Y(_03707_));
 sky130_fd_sc_hd__o22ai_1 _27719_ (.A1(_03470_),
    .A2(_03692_),
    .B1(_03697_),
    .B2(_03700_),
    .Y(_03708_));
 sky130_fd_sc_hd__o211ai_2 _27720_ (.A1(net181),
    .A2(net179),
    .B1(_03707_),
    .C1(_03708_),
    .Y(_03710_));
 sky130_fd_sc_hd__o21ai_4 _27721_ (.A1(net159),
    .A2(_03691_),
    .B1(_03705_),
    .Y(_03711_));
 sky130_fd_sc_hd__o211ai_4 _27722_ (.A1(_03691_),
    .A2(net159),
    .B1(net176),
    .C1(_03705_),
    .Y(_03712_));
 sky130_fd_sc_hd__and3_1 _27723_ (.A(_03710_),
    .B(net178),
    .C(_03706_),
    .X(_03713_));
 sky130_fd_sc_hd__nand3_4 _27724_ (.A(_03710_),
    .B(net178),
    .C(_03706_),
    .Y(_03714_));
 sky130_fd_sc_hd__nand2_1 _27725_ (.A(_03712_),
    .B(_03714_),
    .Y(_03715_));
 sky130_fd_sc_hd__o2bb2ai_1 _27726_ (.A1_N(_03493_),
    .A2_N(_03494_),
    .B1(net201),
    .B2(_03483_),
    .Y(_03716_));
 sky130_fd_sc_hd__a31oi_2 _27727_ (.A1(_03486_),
    .A2(_03493_),
    .A3(_03494_),
    .B1(_03484_),
    .Y(_03717_));
 sky130_fd_sc_hd__a22oi_4 _27728_ (.A1(_03712_),
    .A2(_03714_),
    .B1(_03716_),
    .B2(_03486_),
    .Y(_03718_));
 sky130_fd_sc_hd__o22ai_4 _27729_ (.A1(net157),
    .A2(_08712_),
    .B1(_03715_),
    .B2(_03717_),
    .Y(_03719_));
 sky130_fd_sc_hd__o22ai_4 _27730_ (.A1(net149),
    .A2(_03711_),
    .B1(_03718_),
    .B2(_03719_),
    .Y(_03721_));
 sky130_fd_sc_hd__inv_2 _27731_ (.A(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__o21ai_2 _27732_ (.A1(_09122_),
    .A2(_09123_),
    .B1(_03721_),
    .Y(_03723_));
 sky130_fd_sc_hd__inv_2 _27733_ (.A(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__o21a_1 _27734_ (.A1(_08307_),
    .A2(net216),
    .B1(_03721_),
    .X(_03725_));
 sky130_fd_sc_hd__o21ai_4 _27735_ (.A1(_08307_),
    .A2(net216),
    .B1(_03721_),
    .Y(_03726_));
 sky130_fd_sc_hd__o221ai_4 _27736_ (.A1(net149),
    .A2(_03711_),
    .B1(_03718_),
    .B2(_03719_),
    .C1(net201),
    .Y(_03727_));
 sky130_fd_sc_hd__o2111ai_4 _27737_ (.A1(_02754_),
    .A2(_02746_),
    .B1(_02753_),
    .C1(_03011_),
    .D1(_03013_),
    .Y(_03728_));
 sky130_fd_sc_hd__a211oi_4 _27738_ (.A1(_03253_),
    .A2(_03275_),
    .B1(_03728_),
    .C1(_03279_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand2_1 _27739_ (.A(_03509_),
    .B(_03729_),
    .Y(_03730_));
 sky130_fd_sc_hd__o211ai_4 _27740_ (.A1(_03516_),
    .A2(_03508_),
    .B1(_03512_),
    .C1(_03730_),
    .Y(_03733_));
 sky130_fd_sc_hd__nand3_2 _27741_ (.A(_03509_),
    .B(_03512_),
    .C(_03729_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand4_4 _27742_ (.A(_02760_),
    .B(_03509_),
    .C(_03512_),
    .D(_03729_),
    .Y(_03735_));
 sky130_fd_sc_hd__o21ai_2 _27743_ (.A1(_02759_),
    .A2(_03734_),
    .B1(_03733_),
    .Y(_03736_));
 sky130_fd_sc_hd__a22oi_2 _27744_ (.A1(_03726_),
    .A2(_03727_),
    .B1(_03733_),
    .B2(_03735_),
    .Y(_03737_));
 sky130_fd_sc_hd__a22o_2 _27745_ (.A1(_03726_),
    .A2(_03727_),
    .B1(_03733_),
    .B2(_03735_),
    .X(_03738_));
 sky130_fd_sc_hd__o21a_1 _27746_ (.A1(net197),
    .A2(_03721_),
    .B1(_03735_),
    .X(_03739_));
 sky130_fd_sc_hd__o211ai_4 _27747_ (.A1(_03734_),
    .A2(_02759_),
    .B1(_03727_),
    .C1(_03733_),
    .Y(_03740_));
 sky130_fd_sc_hd__o2111a_1 _27748_ (.A1(net197),
    .A2(_03721_),
    .B1(_03726_),
    .C1(_03733_),
    .D1(_03735_),
    .X(_03741_));
 sky130_fd_sc_hd__o2111ai_4 _27749_ (.A1(net197),
    .A2(_03721_),
    .B1(_03726_),
    .C1(_03733_),
    .D1(_03735_),
    .Y(_03742_));
 sky130_fd_sc_hd__a311oi_2 _27750_ (.A1(_03726_),
    .A2(_03739_),
    .A3(_03733_),
    .B1(_09124_),
    .C1(_03737_),
    .Y(_03744_));
 sky130_fd_sc_hd__o221ai_4 _27751_ (.A1(net148),
    .A2(net147),
    .B1(_03725_),
    .B2(_03740_),
    .C1(_03738_),
    .Y(_03745_));
 sky130_fd_sc_hd__a31oi_4 _27752_ (.A1(net145),
    .A2(_03738_),
    .A3(_03742_),
    .B1(_03724_),
    .Y(_03746_));
 sky130_fd_sc_hd__a2bb2o_2 _27753_ (.A1_N(_09559_),
    .A2_N(_09560_),
    .B1(_03723_),
    .B2(_03745_),
    .X(_03747_));
 sky130_fd_sc_hd__inv_2 _27754_ (.A(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__o311a_2 _27755_ (.A1(_09124_),
    .A2(_03737_),
    .A3(_03741_),
    .B1(_03723_),
    .C1(_07935_),
    .X(_03749_));
 sky130_fd_sc_hd__a311o_2 _27756_ (.A1(net145),
    .A2(_03738_),
    .A3(_03742_),
    .B1(_03724_),
    .C1(_07936_),
    .X(_03750_));
 sky130_fd_sc_hd__a21oi_1 _27757_ (.A1(_03723_),
    .A2(_03745_),
    .B1(_07935_),
    .Y(_03751_));
 sky130_fd_sc_hd__o22ai_4 _27758_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_03724_),
    .B2(_03744_),
    .Y(_03752_));
 sky130_fd_sc_hd__a31o_1 _27759_ (.A1(_03292_),
    .A2(_03527_),
    .A3(_03532_),
    .B1(_03534_),
    .X(_03753_));
 sky130_fd_sc_hd__a21oi_2 _27760_ (.A1(_03528_),
    .A2(_03532_),
    .B1(_03534_),
    .Y(_03755_));
 sky130_fd_sc_hd__a21oi_2 _27761_ (.A1(_03750_),
    .A2(_03752_),
    .B1(_03753_),
    .Y(_03756_));
 sky130_fd_sc_hd__o21ai_1 _27762_ (.A1(_03749_),
    .A2(_03751_),
    .B1(_03755_),
    .Y(_03757_));
 sky130_fd_sc_hd__o21ai_2 _27763_ (.A1(_07935_),
    .A2(_03746_),
    .B1(_03753_),
    .Y(_03758_));
 sky130_fd_sc_hd__a31oi_1 _27764_ (.A1(_03750_),
    .A2(_03752_),
    .A3(_03753_),
    .B1(_09562_),
    .Y(_03759_));
 sky130_fd_sc_hd__o22ai_4 _27765_ (.A1(net156),
    .A2(net154),
    .B1(_03749_),
    .B2(_03758_),
    .Y(_03760_));
 sky130_fd_sc_hd__o211ai_2 _27766_ (.A1(_03758_),
    .A2(_03749_),
    .B1(net144),
    .C1(_03757_),
    .Y(_03761_));
 sky130_fd_sc_hd__o22ai_4 _27767_ (.A1(net144),
    .A2(_03746_),
    .B1(_03756_),
    .B2(_03760_),
    .Y(_03762_));
 sky130_fd_sc_hd__or3_1 _27768_ (.A(net142),
    .B(_09573_),
    .C(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__nand2_1 _27769_ (.A(_03545_),
    .B(_03550_),
    .Y(_03764_));
 sky130_fd_sc_hd__a32o_1 _27770_ (.A1(_07246_),
    .A2(_03539_),
    .A3(_03542_),
    .B1(_03307_),
    .B2(_03326_),
    .X(_03766_));
 sky130_fd_sc_hd__o21ai_1 _27771_ (.A1(_03546_),
    .A2(_03550_),
    .B1(_03545_),
    .Y(_03767_));
 sky130_fd_sc_hd__a31o_1 _27772_ (.A1(_03307_),
    .A2(_03326_),
    .A3(_03545_),
    .B1(_03546_),
    .X(_03768_));
 sky130_fd_sc_hd__a211oi_2 _27773_ (.A1(_03759_),
    .A2(_03757_),
    .B1(_03748_),
    .C1(_07565_),
    .Y(_03769_));
 sky130_fd_sc_hd__o221ai_4 _27774_ (.A1(net144),
    .A2(_03746_),
    .B1(_03756_),
    .B2(_03760_),
    .C1(_07564_),
    .Y(_03770_));
 sky130_fd_sc_hd__a22oi_4 _27775_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_03747_),
    .B2(_03761_),
    .Y(_03771_));
 sky130_fd_sc_hd__o21ai_1 _27776_ (.A1(net221),
    .A2(net219),
    .B1(_03762_),
    .Y(_03772_));
 sky130_fd_sc_hd__nand3_1 _27777_ (.A(_03768_),
    .B(_03770_),
    .C(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__o2bb2ai_1 _27778_ (.A1_N(_03545_),
    .A2_N(_03766_),
    .B1(_03769_),
    .B2(_03771_),
    .Y(_03774_));
 sky130_fd_sc_hd__o211ai_2 _27779_ (.A1(net142),
    .A2(_09573_),
    .B1(_03773_),
    .C1(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__a22o_1 _27780_ (.A1(_09575_),
    .A2(_09577_),
    .B1(_03747_),
    .B2(_03761_),
    .X(_03777_));
 sky130_fd_sc_hd__o2111ai_1 _27781_ (.A1(_07247_),
    .A2(_03543_),
    .B1(_03764_),
    .C1(_03770_),
    .D1(_03772_),
    .Y(_03778_));
 sky130_fd_sc_hd__o2bb2ai_1 _27782_ (.A1_N(_03547_),
    .A2_N(_03764_),
    .B1(_03769_),
    .B2(_03771_),
    .Y(_03779_));
 sky130_fd_sc_hd__o211ai_1 _27783_ (.A1(net142),
    .A2(_09573_),
    .B1(_03778_),
    .C1(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__o21ai_1 _27784_ (.A1(net132),
    .A2(_03762_),
    .B1(_03775_),
    .Y(_03781_));
 sky130_fd_sc_hd__inv_2 _27785_ (.A(_03781_),
    .Y(_03782_));
 sky130_fd_sc_hd__o211ai_4 _27786_ (.A1(_07242_),
    .A2(net248),
    .B1(_03763_),
    .C1(_03775_),
    .Y(_03783_));
 sky130_fd_sc_hd__and3_1 _27787_ (.A(_03780_),
    .B(_07246_),
    .C(_03777_),
    .X(_03784_));
 sky130_fd_sc_hd__nand3_2 _27788_ (.A(_03780_),
    .B(_07246_),
    .C(_03777_),
    .Y(_03785_));
 sky130_fd_sc_hd__nand2_1 _27789_ (.A(_03783_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__a22oi_1 _27790_ (.A1(net226),
    .A2(_03558_),
    .B1(_03572_),
    .B2(_03574_),
    .Y(_03788_));
 sky130_fd_sc_hd__o2bb2ai_1 _27791_ (.A1_N(_03572_),
    .A2_N(_03574_),
    .B1(_06922_),
    .B2(_03559_),
    .Y(_03789_));
 sky130_fd_sc_hd__o22ai_1 _27792_ (.A1(_06922_),
    .A2(_03559_),
    .B1(_03571_),
    .B2(_03584_),
    .Y(_03790_));
 sky130_fd_sc_hd__and4_1 _27793_ (.A(_03560_),
    .B(_03585_),
    .C(_03783_),
    .D(_03785_),
    .X(_03791_));
 sky130_fd_sc_hd__o2bb2ai_2 _27794_ (.A1_N(_03790_),
    .A2_N(_03786_),
    .B1(net140),
    .B2(net141),
    .Y(_03792_));
 sky130_fd_sc_hd__or3_1 _27795_ (.A(net141),
    .B(net140),
    .C(_03781_),
    .X(_03793_));
 sky130_fd_sc_hd__o21ai_1 _27796_ (.A1(_03562_),
    .A2(_03788_),
    .B1(_03786_),
    .Y(_03794_));
 sky130_fd_sc_hd__o2111ai_4 _27797_ (.A1(net226),
    .A2(_03558_),
    .B1(_03783_),
    .C1(_03785_),
    .D1(_03789_),
    .Y(_03795_));
 sky130_fd_sc_hd__nand3_1 _27798_ (.A(net130),
    .B(_03794_),
    .C(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__o22a_2 _27799_ (.A1(net131),
    .A2(_03782_),
    .B1(_03791_),
    .B2(_03792_),
    .X(_03797_));
 sky130_fd_sc_hd__inv_2 _27800_ (.A(_03797_),
    .Y(_03799_));
 sky130_fd_sc_hd__o221a_1 _27801_ (.A1(net130),
    .A2(_03782_),
    .B1(_03791_),
    .B2(_03792_),
    .C1(net226),
    .X(_03800_));
 sky130_fd_sc_hd__o221ai_4 _27802_ (.A1(net131),
    .A2(_03782_),
    .B1(_03791_),
    .B2(_03792_),
    .C1(net226),
    .Y(_03801_));
 sky130_fd_sc_hd__nand3_1 _27803_ (.A(_03796_),
    .B(_06922_),
    .C(_03793_),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_1 _27804_ (.A(_03801_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__nand4_1 _27805_ (.A(_02820_),
    .B(_02822_),
    .C(_03082_),
    .D(_03083_),
    .Y(_03804_));
 sky130_fd_sc_hd__a21oi_1 _27806_ (.A1(_03350_),
    .A2(_06315_),
    .B1(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__nor3_1 _27807_ (.A(_03352_),
    .B(_03804_),
    .C(_03354_),
    .Y(_03806_));
 sky130_fd_sc_hd__o211ai_2 _27808_ (.A1(_06315_),
    .A2(_03350_),
    .B1(_03805_),
    .C1(_03592_),
    .Y(_03807_));
 sky130_fd_sc_hd__o211ai_4 _27809_ (.A1(_03598_),
    .A2(_03591_),
    .B1(_03594_),
    .C1(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand4_4 _27810_ (.A(_03806_),
    .B(_03594_),
    .C(_03592_),
    .D(_02830_),
    .Y(_03810_));
 sky130_fd_sc_hd__nand2_1 _27811_ (.A(_03808_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__a21oi_2 _27812_ (.A1(_03808_),
    .A2(_03810_),
    .B1(_03803_),
    .Y(_03812_));
 sky130_fd_sc_hd__a31o_1 _27813_ (.A1(_03803_),
    .A2(_03808_),
    .A3(_03810_),
    .B1(_10953_),
    .X(_03813_));
 sky130_fd_sc_hd__a211o_1 _27814_ (.A1(_03793_),
    .A2(_03796_),
    .B1(net137),
    .C1(net135),
    .X(_03814_));
 sky130_fd_sc_hd__a22o_1 _27815_ (.A1(_03801_),
    .A2(_03802_),
    .B1(_03808_),
    .B2(_03810_),
    .X(_03815_));
 sky130_fd_sc_hd__o211ai_4 _27816_ (.A1(_03797_),
    .A2(net226),
    .B1(_03810_),
    .C1(_03808_),
    .Y(_03816_));
 sky130_fd_sc_hd__o221ai_4 _27817_ (.A1(net137),
    .A2(net135),
    .B1(_03800_),
    .B2(_03816_),
    .C1(_03815_),
    .Y(_03817_));
 sky130_fd_sc_hd__o31a_1 _27818_ (.A1(net137),
    .A2(net135),
    .A3(_03799_),
    .B1(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__nand3_2 _27819_ (.A(_03817_),
    .B(_06629_),
    .C(_03814_),
    .Y(_03819_));
 sky130_fd_sc_hd__o221a_1 _27820_ (.A1(_10954_),
    .A2(_03797_),
    .B1(_03812_),
    .B2(_03813_),
    .C1(_06630_),
    .X(_03821_));
 sky130_fd_sc_hd__o221ai_4 _27821_ (.A1(_10954_),
    .A2(_03797_),
    .B1(_03812_),
    .B2(_03813_),
    .C1(_06630_),
    .Y(_03822_));
 sky130_fd_sc_hd__o211ai_1 _27822_ (.A1(_06014_),
    .A2(_03363_),
    .B1(_03607_),
    .C1(_03608_),
    .Y(_03823_));
 sky130_fd_sc_hd__o21ai_2 _27823_ (.A1(_06314_),
    .A2(_03605_),
    .B1(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__a21oi_2 _27824_ (.A1(_03819_),
    .A2(_03822_),
    .B1(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__nand3_1 _27825_ (.A(_03819_),
    .B(_03822_),
    .C(_03824_),
    .Y(_03826_));
 sky130_fd_sc_hd__a31o_1 _27826_ (.A1(_03819_),
    .A2(_03822_),
    .A3(_03824_),
    .B1(_11464_),
    .X(_03827_));
 sky130_fd_sc_hd__o22ai_1 _27827_ (.A1(_11465_),
    .A2(_03818_),
    .B1(_03825_),
    .B2(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__o21ai_1 _27828_ (.A1(net284),
    .A2(net281),
    .B1(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__o221ai_4 _27829_ (.A1(_11465_),
    .A2(_03818_),
    .B1(_03825_),
    .B2(_03827_),
    .C1(_06314_),
    .Y(_03830_));
 sky130_fd_sc_hd__a32oi_2 _27830_ (.A1(_03383_),
    .A2(_03618_),
    .A3(_03620_),
    .B1(_03614_),
    .B2(_03616_),
    .Y(_03832_));
 sky130_fd_sc_hd__a21oi_1 _27831_ (.A1(_03829_),
    .A2(_03830_),
    .B1(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__o21bai_2 _27832_ (.A1(_11944_),
    .A2(_03833_),
    .B1_N(_03828_),
    .Y(_03834_));
 sky130_fd_sc_hd__a21oi_1 _27833_ (.A1(_05119_),
    .A2(_03627_),
    .B1(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__o311a_1 _27834_ (.A1(_03615_),
    .A2(_03623_),
    .A3(_03387_),
    .B1(_03834_),
    .C1(_05119_),
    .X(_03836_));
 sky130_fd_sc_hd__nor2_1 _27835_ (.A(_03835_),
    .B(_03836_),
    .Y(net108));
 sky130_fd_sc_hd__or4_2 _27836_ (.A(_03615_),
    .B(_03623_),
    .C(_03834_),
    .D(_03387_),
    .X(_03837_));
 sky130_fd_sc_hd__o2111a_1 _27837_ (.A1(_03630_),
    .A2(_10970_),
    .B1(_06903_),
    .C1(_11471_),
    .D1(_03640_),
    .X(_03838_));
 sky130_fd_sc_hd__a31o_1 _27838_ (.A1(_11471_),
    .A2(_03634_),
    .A3(_03640_),
    .B1(_06904_),
    .X(_03839_));
 sky130_fd_sc_hd__o311a_1 _27839_ (.A1(_11470_),
    .A2(_03633_),
    .A3(_03639_),
    .B1(_07232_),
    .C1(_06903_),
    .X(_03840_));
 sky130_fd_sc_hd__or4_1 _27840_ (.A(_06904_),
    .B(net207),
    .C(net204),
    .D(_03838_),
    .X(_03843_));
 sky130_fd_sc_hd__o311a_1 _27841_ (.A1(_11470_),
    .A2(_03633_),
    .A3(_03639_),
    .B1(_10971_),
    .C1(_06903_),
    .X(_03844_));
 sky130_fd_sc_hd__or4_1 _27842_ (.A(_06897_),
    .B(_06898_),
    .C(_10970_),
    .D(_03838_),
    .X(_03845_));
 sky130_fd_sc_hd__o22a_1 _27843_ (.A1(_10965_),
    .A2(_10967_),
    .B1(_06904_),
    .B2(_03838_),
    .X(_03846_));
 sky130_fd_sc_hd__nor2_2 _27844_ (.A(_03844_),
    .B(_03846_),
    .Y(_03847_));
 sky130_fd_sc_hd__o21ai_2 _27845_ (.A1(_03648_),
    .A2(_03652_),
    .B1(_03647_),
    .Y(_03848_));
 sky130_fd_sc_hd__nand2_2 _27846_ (.A(_03848_),
    .B(_03847_),
    .Y(_03849_));
 sky130_fd_sc_hd__o221ai_4 _27847_ (.A1(net207),
    .A2(net204),
    .B1(_03847_),
    .B2(_03848_),
    .C1(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__o21ai_4 _27848_ (.A1(_07233_),
    .A2(_03839_),
    .B1(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__a21oi_1 _27849_ (.A1(_03843_),
    .A2(_03850_),
    .B1(net150),
    .Y(_03852_));
 sky130_fd_sc_hd__o21ai_4 _27850_ (.A1(_10487_),
    .A2(net165),
    .B1(_03851_),
    .Y(_03854_));
 sky130_fd_sc_hd__o21ai_2 _27851_ (.A1(net164),
    .A2(_10490_),
    .B1(_03850_),
    .Y(_03855_));
 sky130_fd_sc_hd__and3_1 _27852_ (.A(_03850_),
    .B(net150),
    .C(_03843_),
    .X(_03856_));
 sky130_fd_sc_hd__a21o_1 _27853_ (.A1(_03668_),
    .A2(_03670_),
    .B1(_03662_),
    .X(_03857_));
 sky130_fd_sc_hd__a31oi_2 _27854_ (.A1(_03664_),
    .A2(_03668_),
    .A3(_03670_),
    .B1(_03662_),
    .Y(_03858_));
 sky130_fd_sc_hd__o2111ai_4 _27855_ (.A1(_03855_),
    .A2(_03840_),
    .B1(_03672_),
    .C1(_03663_),
    .D1(_03854_),
    .Y(_03859_));
 sky130_fd_sc_hd__o211ai_2 _27856_ (.A1(_03852_),
    .A2(_03856_),
    .B1(_03857_),
    .C1(_03664_),
    .Y(_03860_));
 sky130_fd_sc_hd__o2111ai_1 _27857_ (.A1(_03855_),
    .A2(_03840_),
    .B1(_03664_),
    .C1(_03854_),
    .D1(_03857_),
    .Y(_03861_));
 sky130_fd_sc_hd__o21ai_1 _27858_ (.A1(_03852_),
    .A2(_03856_),
    .B1(_03858_),
    .Y(_03862_));
 sky130_fd_sc_hd__o211ai_4 _27859_ (.A1(_07544_),
    .A2(_07546_),
    .B1(_03859_),
    .C1(_03860_),
    .Y(_03863_));
 sky130_fd_sc_hd__a211o_1 _27860_ (.A1(_03843_),
    .A2(_03850_),
    .B1(_07544_),
    .C1(_07546_),
    .X(_03865_));
 sky130_fd_sc_hd__nand3_1 _27861_ (.A(_03861_),
    .B(_03862_),
    .C(_07548_),
    .Y(_03866_));
 sky130_fd_sc_hd__o21ai_2 _27862_ (.A1(_07548_),
    .A2(_03851_),
    .B1(_03863_),
    .Y(_03867_));
 sky130_fd_sc_hd__o311a_1 _27863_ (.A1(_07544_),
    .A2(_03851_),
    .A3(_07546_),
    .B1(net151),
    .C1(_03863_),
    .X(_03868_));
 sky130_fd_sc_hd__o211ai_4 _27864_ (.A1(_03851_),
    .A2(_07548_),
    .B1(net151),
    .C1(_03863_),
    .Y(_03869_));
 sky130_fd_sc_hd__o211ai_4 _27865_ (.A1(net167),
    .A2(_10024_),
    .B1(_03865_),
    .C1(_03866_),
    .Y(_03870_));
 sky130_fd_sc_hd__nand2_1 _27866_ (.A(_03869_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__and4_1 _27867_ (.A(_02967_),
    .B(_02969_),
    .C(_03220_),
    .D(_03222_),
    .X(_03872_));
 sky130_fd_sc_hd__nand3_1 _27868_ (.A(_03681_),
    .B(_03872_),
    .C(_03456_),
    .Y(_03873_));
 sky130_fd_sc_hd__o211ai_4 _27869_ (.A1(_03685_),
    .A2(_03680_),
    .B1(_03683_),
    .C1(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__nor4b_1 _27870_ (.A(_02866_),
    .B(_03452_),
    .C(_03453_),
    .D_N(_03872_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand3_4 _27871_ (.A(_03876_),
    .B(_03683_),
    .C(_03681_),
    .Y(_03877_));
 sky130_fd_sc_hd__nand3_1 _27872_ (.A(_03871_),
    .B(_03874_),
    .C(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__a21o_1 _27873_ (.A1(_03874_),
    .A2(_03877_),
    .B1(_03871_),
    .X(_03879_));
 sky130_fd_sc_hd__a22o_1 _27874_ (.A1(_03869_),
    .A2(_03870_),
    .B1(_03874_),
    .B2(_03877_),
    .X(_03880_));
 sky130_fd_sc_hd__nand3_1 _27875_ (.A(_03870_),
    .B(_03874_),
    .C(_03877_),
    .Y(_03881_));
 sky130_fd_sc_hd__nand4_2 _27876_ (.A(_03869_),
    .B(_03870_),
    .C(_03874_),
    .D(_03877_),
    .Y(_03882_));
 sky130_fd_sc_hd__nand3_2 _27877_ (.A(_03880_),
    .B(_03882_),
    .C(_07916_),
    .Y(_03883_));
 sky130_fd_sc_hd__o311a_1 _27878_ (.A1(_07544_),
    .A2(_03851_),
    .A3(_07546_),
    .B1(_07917_),
    .C1(_03863_),
    .X(_03884_));
 sky130_fd_sc_hd__or3_1 _27879_ (.A(net183),
    .B(net182),
    .C(_03867_),
    .X(_03885_));
 sky130_fd_sc_hd__o21ai_2 _27880_ (.A1(_07909_),
    .A2(_07911_),
    .B1(_03867_),
    .Y(_03887_));
 sky130_fd_sc_hd__o211ai_2 _27881_ (.A1(net183),
    .A2(net182),
    .B1(_03878_),
    .C1(_03879_),
    .Y(_03888_));
 sky130_fd_sc_hd__and3_2 _27882_ (.A(_08301_),
    .B(_03887_),
    .C(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__a211o_1 _27883_ (.A1(_03883_),
    .A2(_03885_),
    .B1(net181),
    .C1(net179),
    .X(_03890_));
 sky130_fd_sc_hd__a311oi_4 _27884_ (.A1(_03880_),
    .A2(_03882_),
    .A3(_07916_),
    .B1(_03884_),
    .C1(net171),
    .Y(_03891_));
 sky130_fd_sc_hd__nand3_4 _27885_ (.A(_03883_),
    .B(_03885_),
    .C(_09594_),
    .Y(_03892_));
 sky130_fd_sc_hd__o211ai_4 _27886_ (.A1(net189),
    .A2(net186),
    .B1(_03887_),
    .C1(_03888_),
    .Y(_03893_));
 sky130_fd_sc_hd__a21oi_1 _27887_ (.A1(_09140_),
    .A2(_03691_),
    .B1(_03695_),
    .Y(_03894_));
 sky130_fd_sc_hd__a31o_1 _27888_ (.A1(_03471_),
    .A2(_03693_),
    .A3(_03699_),
    .B1(_03700_),
    .X(_03895_));
 sky130_fd_sc_hd__a21oi_1 _27889_ (.A1(_03695_),
    .A2(_03699_),
    .B1(_03700_),
    .Y(_03896_));
 sky130_fd_sc_hd__o2bb2ai_4 _27890_ (.A1_N(_03892_),
    .A2_N(_03893_),
    .B1(_03894_),
    .B2(_03697_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand3_2 _27891_ (.A(_03895_),
    .B(_03893_),
    .C(_03892_),
    .Y(_03899_));
 sky130_fd_sc_hd__nand3_1 _27892_ (.A(_03898_),
    .B(_03899_),
    .C(net159),
    .Y(_03900_));
 sky130_fd_sc_hd__a31o_2 _27893_ (.A1(_03898_),
    .A2(_03899_),
    .A3(net159),
    .B1(_03889_),
    .X(_03901_));
 sky130_fd_sc_hd__o311a_1 _27894_ (.A1(_08311_),
    .A2(_03483_),
    .A3(net215),
    .B1(_03712_),
    .C1(_03502_),
    .X(_03902_));
 sky130_fd_sc_hd__o221ai_4 _27895_ (.A1(net201),
    .A2(_03483_),
    .B1(net178),
    .B2(_03711_),
    .C1(_03502_),
    .Y(_03903_));
 sky130_fd_sc_hd__a31oi_2 _27896_ (.A1(_03485_),
    .A2(_03502_),
    .A3(_03712_),
    .B1(_03713_),
    .Y(_03904_));
 sky130_fd_sc_hd__a31oi_1 _27897_ (.A1(_03898_),
    .A2(_03899_),
    .A3(net159),
    .B1(_09140_),
    .Y(_03905_));
 sky130_fd_sc_hd__a311oi_4 _27898_ (.A1(_03898_),
    .A2(_03899_),
    .A3(net159),
    .B1(_09140_),
    .C1(_03889_),
    .Y(_03906_));
 sky130_fd_sc_hd__a311o_1 _27899_ (.A1(_03898_),
    .A2(_03899_),
    .A3(net159),
    .B1(_09140_),
    .C1(_03889_),
    .X(_03907_));
 sky130_fd_sc_hd__a2bb2oi_2 _27900_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_03890_),
    .B2(_03900_),
    .Y(_03909_));
 sky130_fd_sc_hd__a2bb2o_1 _27901_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_03890_),
    .B2(_03900_),
    .X(_03910_));
 sky130_fd_sc_hd__o211ai_1 _27902_ (.A1(_03713_),
    .A2(_03902_),
    .B1(_03907_),
    .C1(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__o21ai_1 _27903_ (.A1(_03906_),
    .A2(_03909_),
    .B1(_03904_),
    .Y(_03912_));
 sky130_fd_sc_hd__nand3_2 _27904_ (.A(_03911_),
    .B(_03912_),
    .C(net149),
    .Y(_03913_));
 sky130_fd_sc_hd__a22o_1 _27905_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_03890_),
    .B2(_03900_),
    .X(_03914_));
 sky130_fd_sc_hd__nand3_1 _27906_ (.A(_03910_),
    .B(_03904_),
    .C(_03907_),
    .Y(_03915_));
 sky130_fd_sc_hd__o2bb2ai_1 _27907_ (.A1_N(_03714_),
    .A2_N(_03903_),
    .B1(_03906_),
    .B2(_03909_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand3_1 _27908_ (.A(_03915_),
    .B(_03916_),
    .C(net149),
    .Y(_03917_));
 sky130_fd_sc_hd__o21ai_4 _27909_ (.A1(net149),
    .A2(_03901_),
    .B1(_03913_),
    .Y(_03918_));
 sky130_fd_sc_hd__o211ai_4 _27910_ (.A1(_03901_),
    .A2(net149),
    .B1(net176),
    .C1(_03913_),
    .Y(_03920_));
 sky130_fd_sc_hd__o211ai_4 _27911_ (.A1(_08728_),
    .A2(_08729_),
    .B1(_03914_),
    .C1(_03917_),
    .Y(_03921_));
 sky130_fd_sc_hd__nand2_2 _27912_ (.A(_03920_),
    .B(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__a31oi_2 _27913_ (.A1(_03727_),
    .A2(_03733_),
    .A3(_03735_),
    .B1(_03725_),
    .Y(_03923_));
 sky130_fd_sc_hd__o311a_2 _27914_ (.A1(_08311_),
    .A2(net215),
    .A3(_03722_),
    .B1(_03740_),
    .C1(_03922_),
    .X(_03924_));
 sky130_fd_sc_hd__a21o_1 _27915_ (.A1(_03726_),
    .A2(_03740_),
    .B1(_03922_),
    .X(_03925_));
 sky130_fd_sc_hd__o21ai_4 _27916_ (.A1(_03922_),
    .A2(_03923_),
    .B1(net145),
    .Y(_03926_));
 sky130_fd_sc_hd__o32a_2 _27917_ (.A1(net148),
    .A2(net147),
    .A3(_03918_),
    .B1(_03924_),
    .B2(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__o22ai_4 _27918_ (.A1(net145),
    .A2(_03918_),
    .B1(_03924_),
    .B2(_03926_),
    .Y(_03928_));
 sky130_fd_sc_hd__and3_1 _27919_ (.A(_09554_),
    .B(_09557_),
    .C(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__or3_4 _27920_ (.A(net156),
    .B(net154),
    .C(_03927_),
    .X(_03931_));
 sky130_fd_sc_hd__o21a_2 _27921_ (.A1(_08307_),
    .A2(net216),
    .B1(_03928_),
    .X(_03932_));
 sky130_fd_sc_hd__o21ai_4 _27922_ (.A1(_08307_),
    .A2(net216),
    .B1(_03928_),
    .Y(_03933_));
 sky130_fd_sc_hd__o221ai_4 _27923_ (.A1(net145),
    .A2(_03918_),
    .B1(_03924_),
    .B2(_03926_),
    .C1(net201),
    .Y(_03934_));
 sky130_fd_sc_hd__nor3_1 _27924_ (.A(_03030_),
    .B(_03291_),
    .C(_03293_),
    .Y(_03935_));
 sky130_fd_sc_hd__o211ai_2 _27925_ (.A1(_03506_),
    .A2(_03530_),
    .B1(_03935_),
    .C1(_03535_),
    .Y(_03936_));
 sky130_fd_sc_hd__a31o_1 _27926_ (.A1(_03745_),
    .A2(_07935_),
    .A3(_03723_),
    .B1(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__o211ai_4 _27927_ (.A1(_03755_),
    .A2(_03749_),
    .B1(_03752_),
    .C1(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__a21oi_2 _27928_ (.A1(_03035_),
    .A2(_03037_),
    .B1(_03936_),
    .Y(_03939_));
 sky130_fd_sc_hd__nand3_4 _27929_ (.A(_03750_),
    .B(_03752_),
    .C(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__nand2_2 _27930_ (.A(_03938_),
    .B(_03940_),
    .Y(_03942_));
 sky130_fd_sc_hd__inv_2 _27931_ (.A(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__a22oi_2 _27932_ (.A1(_03933_),
    .A2(_03934_),
    .B1(_03938_),
    .B2(_03940_),
    .Y(_03944_));
 sky130_fd_sc_hd__a22o_1 _27933_ (.A1(_03933_),
    .A2(_03934_),
    .B1(_03938_),
    .B2(_03940_),
    .X(_03945_));
 sky130_fd_sc_hd__o211ai_4 _27934_ (.A1(net197),
    .A2(_03928_),
    .B1(_03938_),
    .C1(_03940_),
    .Y(_03946_));
 sky130_fd_sc_hd__o2111a_1 _27935_ (.A1(net197),
    .A2(_03928_),
    .B1(_03933_),
    .C1(_03938_),
    .D1(_03940_),
    .X(_03947_));
 sky130_fd_sc_hd__o2111ai_1 _27936_ (.A1(net197),
    .A2(_03928_),
    .B1(_03933_),
    .C1(_03938_),
    .D1(_03940_),
    .Y(_03948_));
 sky130_fd_sc_hd__nor3b_1 _27937_ (.A(_09562_),
    .B(_03944_),
    .C_N(_03948_),
    .Y(_03949_));
 sky130_fd_sc_hd__o221ai_4 _27938_ (.A1(net156),
    .A2(net154),
    .B1(_03932_),
    .B2(_03946_),
    .C1(_03945_),
    .Y(_03950_));
 sky130_fd_sc_hd__a22o_4 _27939_ (.A1(_09575_),
    .A2(_09577_),
    .B1(_03931_),
    .B2(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__inv_2 _27940_ (.A(_03951_),
    .Y(_03954_));
 sky130_fd_sc_hd__o311a_4 _27941_ (.A1(_09562_),
    .A2(_03944_),
    .A3(_03947_),
    .B1(_03931_),
    .C1(_07935_),
    .X(_03955_));
 sky130_fd_sc_hd__nand3_4 _27942_ (.A(_03950_),
    .B(_07935_),
    .C(_03931_),
    .Y(_03956_));
 sky130_fd_sc_hd__a21oi_4 _27943_ (.A1(_03931_),
    .A2(_03950_),
    .B1(_07935_),
    .Y(_03957_));
 sky130_fd_sc_hd__o22ai_4 _27944_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_03929_),
    .B2(_03949_),
    .Y(_03958_));
 sky130_fd_sc_hd__a31o_1 _27945_ (.A1(_03547_),
    .A2(_03764_),
    .A3(_03770_),
    .B1(_03771_),
    .X(_03959_));
 sky130_fd_sc_hd__a21oi_4 _27946_ (.A1(_03767_),
    .A2(_03770_),
    .B1(_03771_),
    .Y(_03960_));
 sky130_fd_sc_hd__o21ai_4 _27947_ (.A1(_03955_),
    .A2(_03957_),
    .B1(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__a31oi_4 _27948_ (.A1(_03956_),
    .A2(_03958_),
    .A3(_03959_),
    .B1(_09578_),
    .Y(_03962_));
 sky130_fd_sc_hd__o311a_2 _27949_ (.A1(_03955_),
    .A2(_03960_),
    .A3(_03957_),
    .B1(net132),
    .C1(_03961_),
    .X(_03963_));
 sky130_fd_sc_hd__o311ai_4 _27950_ (.A1(_03955_),
    .A2(_03960_),
    .A3(_03957_),
    .B1(net132),
    .C1(_03961_),
    .Y(_03965_));
 sky130_fd_sc_hd__a21oi_1 _27951_ (.A1(_03962_),
    .A2(_03961_),
    .B1(_03954_),
    .Y(_03966_));
 sky130_fd_sc_hd__o311a_1 _27952_ (.A1(_06918_),
    .A2(_03559_),
    .A3(net249),
    .B1(_03783_),
    .C1(_03585_),
    .X(_03967_));
 sky130_fd_sc_hd__a31oi_4 _27953_ (.A1(_03560_),
    .A2(_03585_),
    .A3(_03783_),
    .B1(_03784_),
    .Y(_03968_));
 sky130_fd_sc_hd__a22oi_4 _27954_ (.A1(_07561_),
    .A2(_07563_),
    .B1(_03962_),
    .B2(_03961_),
    .Y(_03969_));
 sky130_fd_sc_hd__a211oi_1 _27955_ (.A1(_03962_),
    .A2(_03961_),
    .B1(_03954_),
    .C1(_07565_),
    .Y(_03970_));
 sky130_fd_sc_hd__o211ai_4 _27956_ (.A1(_07560_),
    .A2(net217),
    .B1(_03951_),
    .C1(_03965_),
    .Y(_03971_));
 sky130_fd_sc_hd__a2bb2oi_4 _27957_ (.A1_N(net221),
    .A2_N(net219),
    .B1(_03951_),
    .B2(_03965_),
    .Y(_03972_));
 sky130_fd_sc_hd__o22ai_2 _27958_ (.A1(net221),
    .A2(net219),
    .B1(_03954_),
    .B2(_03963_),
    .Y(_03973_));
 sky130_fd_sc_hd__a21oi_1 _27959_ (.A1(_03951_),
    .A2(_03969_),
    .B1(_03972_),
    .Y(_03974_));
 sky130_fd_sc_hd__o211ai_1 _27960_ (.A1(_03784_),
    .A2(_03967_),
    .B1(_03971_),
    .C1(_03973_),
    .Y(_03976_));
 sky130_fd_sc_hd__o21ai_1 _27961_ (.A1(_03970_),
    .A2(_03972_),
    .B1(_03968_),
    .Y(_03977_));
 sky130_fd_sc_hd__nand3_1 _27962_ (.A(_03973_),
    .B(_03968_),
    .C(_03971_),
    .Y(_03978_));
 sky130_fd_sc_hd__o22ai_2 _27963_ (.A1(_03784_),
    .A2(_03967_),
    .B1(_03970_),
    .B2(_03972_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand3_1 _27964_ (.A(net130),
    .B(_03976_),
    .C(_03977_),
    .Y(_03980_));
 sky130_fd_sc_hd__or3_2 _27965_ (.A(net141),
    .B(net140),
    .C(_03966_),
    .X(_03981_));
 sky130_fd_sc_hd__o211ai_2 _27966_ (.A1(net141),
    .A2(net140),
    .B1(_03978_),
    .C1(_03979_),
    .Y(_03982_));
 sky130_fd_sc_hd__o31a_1 _27967_ (.A1(net130),
    .A2(_03954_),
    .A3(_03963_),
    .B1(_03980_),
    .X(_03983_));
 sky130_fd_sc_hd__o31a_2 _27968_ (.A1(net141),
    .A2(net140),
    .A3(_03966_),
    .B1(_03982_),
    .X(_03984_));
 sky130_fd_sc_hd__a31oi_2 _27969_ (.A1(net130),
    .A2(_03978_),
    .A3(_03979_),
    .B1(_07247_),
    .Y(_03985_));
 sky130_fd_sc_hd__and3_2 _27970_ (.A(_03982_),
    .B(_07246_),
    .C(_03981_),
    .X(_03987_));
 sky130_fd_sc_hd__o21ai_2 _27971_ (.A1(net130),
    .A2(_03966_),
    .B1(_03985_),
    .Y(_03988_));
 sky130_fd_sc_hd__a2bb2oi_2 _27972_ (.A1_N(_07242_),
    .A2_N(net248),
    .B1(_03981_),
    .B2(_03982_),
    .Y(_03989_));
 sky130_fd_sc_hd__o311ai_4 _27973_ (.A1(net130),
    .A2(_03954_),
    .A3(_03963_),
    .B1(_03980_),
    .C1(_07247_),
    .Y(_03990_));
 sky130_fd_sc_hd__o2bb2ai_1 _27974_ (.A1_N(_03801_),
    .A2_N(_03816_),
    .B1(_07246_),
    .B2(_03984_),
    .Y(_03991_));
 sky130_fd_sc_hd__o221ai_4 _27975_ (.A1(_03799_),
    .A2(_06922_),
    .B1(_03989_),
    .B2(_03987_),
    .C1(_03816_),
    .Y(_03992_));
 sky130_fd_sc_hd__o221ai_4 _27976_ (.A1(net137),
    .A2(net135),
    .B1(_03987_),
    .B2(_03991_),
    .C1(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__or3_2 _27977_ (.A(net137),
    .B(net135),
    .C(_03984_),
    .X(_03994_));
 sky130_fd_sc_hd__inv_2 _27978_ (.A(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__a211o_2 _27979_ (.A1(_03993_),
    .A2(_03994_),
    .B1(_11459_),
    .C1(net129),
    .X(_03996_));
 sky130_fd_sc_hd__a21oi_2 _27980_ (.A1(_03993_),
    .A2(_03994_),
    .B1(_06922_),
    .Y(_03998_));
 sky130_fd_sc_hd__a22o_1 _27981_ (.A1(_06915_),
    .A2(_06917_),
    .B1(_03993_),
    .B2(_03994_),
    .X(_03999_));
 sky130_fd_sc_hd__o21ai_1 _27982_ (.A1(_06918_),
    .A2(net249),
    .B1(_03993_),
    .Y(_04000_));
 sky130_fd_sc_hd__o221a_1 _27983_ (.A1(_06918_),
    .A2(net249),
    .B1(_10954_),
    .B2(_03984_),
    .C1(_03993_),
    .X(_04001_));
 sky130_fd_sc_hd__o221ai_4 _27984_ (.A1(_06918_),
    .A2(net249),
    .B1(_10954_),
    .B2(_03984_),
    .C1(_03993_),
    .Y(_04002_));
 sky130_fd_sc_hd__nand4_2 _27985_ (.A(_03609_),
    .B(_03370_),
    .C(_03095_),
    .D(_03608_),
    .Y(_04003_));
 sky130_fd_sc_hd__a31oi_2 _27986_ (.A1(_03817_),
    .A2(_06629_),
    .A3(_03814_),
    .B1(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__a31o_1 _27987_ (.A1(_03817_),
    .A2(_06629_),
    .A3(_03814_),
    .B1(_04003_),
    .X(_04005_));
 sky130_fd_sc_hd__a211oi_1 _27988_ (.A1(_03824_),
    .A2(_03819_),
    .B1(_03821_),
    .C1(_04004_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand3_1 _27989_ (.A(_03822_),
    .B(_03826_),
    .C(_04005_),
    .Y(_04007_));
 sky130_fd_sc_hd__nand3b_1 _27990_ (.A_N(_04003_),
    .B(_03822_),
    .C(_03819_),
    .Y(_04009_));
 sky130_fd_sc_hd__and3_1 _27991_ (.A(_04004_),
    .B(_03822_),
    .C(_03104_),
    .X(_04010_));
 sky130_fd_sc_hd__a31o_1 _27992_ (.A1(_03104_),
    .A2(_03822_),
    .A3(_04004_),
    .B1(_04006_),
    .X(_04011_));
 sky130_fd_sc_hd__o22ai_2 _27993_ (.A1(_03998_),
    .A2(_04001_),
    .B1(_04006_),
    .B2(_04010_),
    .Y(_04012_));
 sky130_fd_sc_hd__o211ai_4 _27994_ (.A1(_04009_),
    .A2(_03103_),
    .B1(_04002_),
    .C1(_04007_),
    .Y(_04013_));
 sky130_fd_sc_hd__o221ai_4 _27995_ (.A1(_11459_),
    .A2(net129),
    .B1(_03998_),
    .B2(_04013_),
    .C1(_04012_),
    .Y(_04014_));
 sky130_fd_sc_hd__and3_1 _27996_ (.A(_04014_),
    .B(_06629_),
    .C(_03996_),
    .X(_04015_));
 sky130_fd_sc_hd__o211ai_2 _27997_ (.A1(_06626_),
    .A2(_06627_),
    .B1(_03996_),
    .C1(_04014_),
    .Y(_04016_));
 sky130_fd_sc_hd__a22o_1 _27998_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_03996_),
    .B2(_04014_),
    .X(_04017_));
 sky130_fd_sc_hd__a21boi_1 _27999_ (.A1(_03832_),
    .A2(_03830_),
    .B1_N(_03829_),
    .Y(_04018_));
 sky130_fd_sc_hd__a21boi_1 _28000_ (.A1(_04016_),
    .A2(_04017_),
    .B1_N(_04018_),
    .Y(_04020_));
 sky130_fd_sc_hd__o211ai_4 _28001_ (.A1(_11944_),
    .A2(_04020_),
    .B1(_04014_),
    .C1(_03996_),
    .Y(_04021_));
 sky130_fd_sc_hd__a21oi_1 _28002_ (.A1(_05119_),
    .A2(_03837_),
    .B1(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__o311a_1 _28003_ (.A1(_03624_),
    .A2(_03834_),
    .A3(_03387_),
    .B1(_04021_),
    .C1(_05119_),
    .X(_04023_));
 sky130_fd_sc_hd__nor2_1 _28004_ (.A(_04022_),
    .B(_04023_),
    .Y(net110));
 sky130_fd_sc_hd__o21ai_1 _28005_ (.A1(_03837_),
    .A2(_04021_),
    .B1(_05119_),
    .Y(_04024_));
 sky130_fd_sc_hd__a211o_1 _28006_ (.A1(_03848_),
    .A2(_03847_),
    .B1(_03844_),
    .C1(_11470_),
    .X(_04025_));
 sky130_fd_sc_hd__a31o_1 _28007_ (.A1(_11471_),
    .A2(_03845_),
    .A3(_03849_),
    .B1(_07232_),
    .X(_04026_));
 sky130_fd_sc_hd__a311o_1 _28008_ (.A1(_11471_),
    .A2(_03845_),
    .A3(_03849_),
    .B1(_07548_),
    .C1(_07232_),
    .X(_04027_));
 sky130_fd_sc_hd__o211a_1 _28009_ (.A1(net207),
    .A2(net204),
    .B1(_10971_),
    .C1(_04025_),
    .X(_04028_));
 sky130_fd_sc_hd__a311o_2 _28010_ (.A1(_11471_),
    .A2(_03845_),
    .A3(_03849_),
    .B1(_10970_),
    .C1(_07232_),
    .X(_04030_));
 sky130_fd_sc_hd__a21oi_1 _28011_ (.A1(_07233_),
    .A2(_04025_),
    .B1(_10971_),
    .Y(_04031_));
 sky130_fd_sc_hd__a22o_1 _28012_ (.A1(_10966_),
    .A2(_10968_),
    .B1(_04025_),
    .B2(_07233_),
    .X(_04032_));
 sky130_fd_sc_hd__o211ai_2 _28013_ (.A1(net152),
    .A2(_03659_),
    .B1(_03672_),
    .C1(_03854_),
    .Y(_04033_));
 sky130_fd_sc_hd__o221ai_4 _28014_ (.A1(_04028_),
    .A2(_04031_),
    .B1(_03856_),
    .B2(_03858_),
    .C1(_03854_),
    .Y(_04034_));
 sky130_fd_sc_hd__o2111ai_4 _28015_ (.A1(_10492_),
    .A2(_03851_),
    .B1(_04030_),
    .C1(_04032_),
    .D1(_04033_),
    .Y(_04035_));
 sky130_fd_sc_hd__nand3_2 _28016_ (.A(_04034_),
    .B(_04035_),
    .C(_07548_),
    .Y(_04036_));
 sky130_fd_sc_hd__and3_1 _28017_ (.A(_07545_),
    .B(_07547_),
    .C(_04026_),
    .X(_04037_));
 sky130_fd_sc_hd__a21oi_2 _28018_ (.A1(_04034_),
    .A2(_04035_),
    .B1(_07550_),
    .Y(_04038_));
 sky130_fd_sc_hd__o21ai_4 _28019_ (.A1(_07548_),
    .A2(_04026_),
    .B1(_04036_),
    .Y(_04039_));
 sky130_fd_sc_hd__a21oi_1 _28020_ (.A1(_04027_),
    .A2(_04036_),
    .B1(net150),
    .Y(_04041_));
 sky130_fd_sc_hd__a2bb2o_1 _28021_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_04027_),
    .B2(_04036_),
    .X(_04042_));
 sky130_fd_sc_hd__and3_1 _28022_ (.A(_04036_),
    .B(net150),
    .C(_04027_),
    .X(_04043_));
 sky130_fd_sc_hd__nor2_1 _28023_ (.A(_04041_),
    .B(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__o2bb2ai_1 _28024_ (.A1_N(_03874_),
    .A2_N(_03877_),
    .B1(net152),
    .B2(_03867_),
    .Y(_04045_));
 sky130_fd_sc_hd__a31oi_2 _28025_ (.A1(_03870_),
    .A2(_03874_),
    .A3(_03877_),
    .B1(_03868_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand3_1 _28026_ (.A(_04044_),
    .B(_03881_),
    .C(_03869_),
    .Y(_04047_));
 sky130_fd_sc_hd__o211ai_1 _28027_ (.A1(_04041_),
    .A2(_04043_),
    .B1(_04045_),
    .C1(_03870_),
    .Y(_04048_));
 sky130_fd_sc_hd__nand3_1 _28028_ (.A(_04044_),
    .B(_04045_),
    .C(_03870_),
    .Y(_04049_));
 sky130_fd_sc_hd__o211ai_1 _28029_ (.A1(_04041_),
    .A2(_04043_),
    .B1(_03869_),
    .C1(_03881_),
    .Y(_04050_));
 sky130_fd_sc_hd__o211ai_2 _28030_ (.A1(net183),
    .A2(net182),
    .B1(_04047_),
    .C1(_04048_),
    .Y(_04052_));
 sky130_fd_sc_hd__nand3_2 _28031_ (.A(_04049_),
    .B(_04050_),
    .C(_07916_),
    .Y(_04053_));
 sky130_fd_sc_hd__o31a_2 _28032_ (.A1(_07916_),
    .A2(_04037_),
    .A3(_04038_),
    .B1(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__o221a_1 _28033_ (.A1(_08293_),
    .A2(_08295_),
    .B1(_04039_),
    .B2(_07916_),
    .C1(_04052_),
    .X(_04055_));
 sky130_fd_sc_hd__inv_2 _28034_ (.A(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__o311a_1 _28035_ (.A1(net183),
    .A2(_04039_),
    .A3(net182),
    .B1(_10027_),
    .C1(_04052_),
    .X(_04057_));
 sky130_fd_sc_hd__o211ai_2 _28036_ (.A1(_04039_),
    .A2(_07916_),
    .B1(_10027_),
    .C1(_04052_),
    .Y(_04058_));
 sky130_fd_sc_hd__o311a_1 _28037_ (.A1(_07916_),
    .A2(_04037_),
    .A3(_04038_),
    .B1(net152),
    .C1(_04053_),
    .X(_04059_));
 sky130_fd_sc_hd__o311ai_4 _28038_ (.A1(_07916_),
    .A2(_04037_),
    .A3(_04038_),
    .B1(net152),
    .C1(_04053_),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2_1 _28039_ (.A(_04058_),
    .B(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__and4_1 _28040_ (.A(_03238_),
    .B(_03240_),
    .C(_03469_),
    .D(_03471_),
    .X(_04064_));
 sky130_fd_sc_hd__nand3_1 _28041_ (.A(_03892_),
    .B(_04064_),
    .C(_03702_),
    .Y(_04065_));
 sky130_fd_sc_hd__o211ai_4 _28042_ (.A1(_03896_),
    .A2(_03891_),
    .B1(_03893_),
    .C1(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__and4_1 _28043_ (.A(_04064_),
    .B(_03701_),
    .C(_03699_),
    .D(_03125_),
    .X(_04067_));
 sky130_fd_sc_hd__nand3_4 _28044_ (.A(_04067_),
    .B(_03893_),
    .C(_03892_),
    .Y(_04068_));
 sky130_fd_sc_hd__nand3_1 _28045_ (.A(_04061_),
    .B(_04066_),
    .C(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__a21o_1 _28046_ (.A1(_04066_),
    .A2(_04068_),
    .B1(_04061_),
    .X(_04070_));
 sky130_fd_sc_hd__a22o_1 _28047_ (.A1(_04058_),
    .A2(_04060_),
    .B1(_04066_),
    .B2(_04068_),
    .X(_04071_));
 sky130_fd_sc_hd__nand3_2 _28048_ (.A(_04060_),
    .B(_04066_),
    .C(_04068_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand4_2 _28049_ (.A(_04058_),
    .B(_04060_),
    .C(_04066_),
    .D(_04068_),
    .Y(_04073_));
 sky130_fd_sc_hd__nand3_2 _28050_ (.A(_04071_),
    .B(_04073_),
    .C(net159),
    .Y(_04075_));
 sky130_fd_sc_hd__o21ai_2 _28051_ (.A1(_08293_),
    .A2(_08295_),
    .B1(_04054_),
    .Y(_04076_));
 sky130_fd_sc_hd__nand3_1 _28052_ (.A(_04070_),
    .B(net159),
    .C(_04069_),
    .Y(_04077_));
 sky130_fd_sc_hd__o31a_1 _28053_ (.A1(net181),
    .A2(net179),
    .A3(_04054_),
    .B1(_04075_),
    .X(_04078_));
 sky130_fd_sc_hd__and3_1 _28054_ (.A(_08715_),
    .B(_04076_),
    .C(_04077_),
    .X(_04079_));
 sky130_fd_sc_hd__a22o_2 _28055_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_04056_),
    .B2(_04075_),
    .X(_04080_));
 sky130_fd_sc_hd__a311oi_2 _28056_ (.A1(_04071_),
    .A2(_04073_),
    .A3(net159),
    .B1(net171),
    .C1(_04055_),
    .Y(_04081_));
 sky130_fd_sc_hd__nand3_4 _28057_ (.A(_04075_),
    .B(_09594_),
    .C(_04056_),
    .Y(_04082_));
 sky130_fd_sc_hd__o211ai_4 _28058_ (.A1(net189),
    .A2(net186),
    .B1(_04076_),
    .C1(_04077_),
    .Y(_04083_));
 sky130_fd_sc_hd__a21oi_1 _28059_ (.A1(_03714_),
    .A2(_03903_),
    .B1(_03909_),
    .Y(_04084_));
 sky130_fd_sc_hd__a31o_1 _28060_ (.A1(_03714_),
    .A2(_03903_),
    .A3(_03907_),
    .B1(_03909_),
    .X(_04086_));
 sky130_fd_sc_hd__a21oi_1 _28061_ (.A1(_03904_),
    .A2(_03907_),
    .B1(_03909_),
    .Y(_04087_));
 sky130_fd_sc_hd__o2bb2ai_2 _28062_ (.A1_N(_04082_),
    .A2_N(_04083_),
    .B1(_04084_),
    .B2(_03906_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand3_2 _28063_ (.A(_04086_),
    .B(_04083_),
    .C(_04082_),
    .Y(_04089_));
 sky130_fd_sc_hd__nand3_2 _28064_ (.A(_04088_),
    .B(_04089_),
    .C(net149),
    .Y(_04090_));
 sky130_fd_sc_hd__a31oi_4 _28065_ (.A1(_04088_),
    .A2(_04089_),
    .A3(net149),
    .B1(_04079_),
    .Y(_04091_));
 sky130_fd_sc_hd__a31o_1 _28066_ (.A1(_04088_),
    .A2(_04089_),
    .A3(net149),
    .B1(_04079_),
    .X(_04092_));
 sky130_fd_sc_hd__o311a_1 _28067_ (.A1(net157),
    .A2(_08712_),
    .A3(_04078_),
    .B1(_09124_),
    .C1(_04090_),
    .X(_04093_));
 sky130_fd_sc_hd__o221ai_4 _28068_ (.A1(net201),
    .A2(_03722_),
    .B1(net178),
    .B2(_03918_),
    .C1(_03740_),
    .Y(_04094_));
 sky130_fd_sc_hd__nand2_1 _28069_ (.A(_03921_),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__a31oi_1 _28070_ (.A1(_04088_),
    .A2(_04089_),
    .A3(net149),
    .B1(_09140_),
    .Y(_04096_));
 sky130_fd_sc_hd__o211a_1 _28071_ (.A1(net149),
    .A2(_04078_),
    .B1(_09139_),
    .C1(_04090_),
    .X(_04097_));
 sky130_fd_sc_hd__nand3_2 _28072_ (.A(_04090_),
    .B(_09139_),
    .C(_04080_),
    .Y(_04098_));
 sky130_fd_sc_hd__a2bb2oi_2 _28073_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_04080_),
    .B2(_04090_),
    .Y(_04099_));
 sky130_fd_sc_hd__a2bb2o_1 _28074_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_04080_),
    .B2(_04090_),
    .X(_04100_));
 sky130_fd_sc_hd__nand3_1 _28075_ (.A(_04095_),
    .B(_04098_),
    .C(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__o2bb2ai_1 _28076_ (.A1_N(_03920_),
    .A2_N(_03925_),
    .B1(_04097_),
    .B2(_04099_),
    .Y(_04102_));
 sky130_fd_sc_hd__o211ai_2 _28077_ (.A1(net148),
    .A2(net147),
    .B1(_04101_),
    .C1(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__o2111ai_4 _28078_ (.A1(_09139_),
    .A2(_04091_),
    .B1(_04094_),
    .C1(_04098_),
    .D1(_03921_),
    .Y(_04104_));
 sky130_fd_sc_hd__o21ai_1 _28079_ (.A1(_04097_),
    .A2(_04099_),
    .B1(_04095_),
    .Y(_04105_));
 sky130_fd_sc_hd__o211ai_4 _28080_ (.A1(net148),
    .A2(net147),
    .B1(_04104_),
    .C1(_04105_),
    .Y(_04107_));
 sky130_fd_sc_hd__o21ai_2 _28081_ (.A1(net145),
    .A2(_04091_),
    .B1(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__a31o_1 _28082_ (.A1(net145),
    .A2(_04101_),
    .A3(_04102_),
    .B1(_04093_),
    .X(_04109_));
 sky130_fd_sc_hd__o211ai_4 _28083_ (.A1(net145),
    .A2(_04092_),
    .B1(_04103_),
    .C1(net176),
    .Y(_04110_));
 sky130_fd_sc_hd__o211a_1 _28084_ (.A1(net145),
    .A2(_04091_),
    .B1(net178),
    .C1(_04107_),
    .X(_04111_));
 sky130_fd_sc_hd__o211ai_4 _28085_ (.A1(net145),
    .A2(_04091_),
    .B1(net178),
    .C1(_04107_),
    .Y(_04112_));
 sky130_fd_sc_hd__nand2_2 _28086_ (.A(_04110_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__a31o_1 _28087_ (.A1(_03934_),
    .A2(_03938_),
    .A3(_03940_),
    .B1(_03932_),
    .X(_04114_));
 sky130_fd_sc_hd__a31oi_4 _28088_ (.A1(_03934_),
    .A2(_03938_),
    .A3(_03940_),
    .B1(_03932_),
    .Y(_04115_));
 sky130_fd_sc_hd__o2111ai_1 _28089_ (.A1(net201),
    .A2(_03927_),
    .B1(_03946_),
    .C1(_04110_),
    .D1(_04112_),
    .Y(_04116_));
 sky130_fd_sc_hd__nand2_1 _28090_ (.A(_04114_),
    .B(_04113_),
    .Y(_04118_));
 sky130_fd_sc_hd__o211ai_2 _28091_ (.A1(net156),
    .A2(net154),
    .B1(_04116_),
    .C1(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__a311o_2 _28092_ (.A1(net145),
    .A2(_04101_),
    .A3(_04102_),
    .B1(net144),
    .C1(_04093_),
    .X(_04120_));
 sky130_fd_sc_hd__o311a_1 _28093_ (.A1(_08311_),
    .A2(net215),
    .A3(_03927_),
    .B1(_03946_),
    .C1(_04113_),
    .X(_04121_));
 sky130_fd_sc_hd__nand2_1 _28094_ (.A(_04113_),
    .B(_04115_),
    .Y(_04122_));
 sky130_fd_sc_hd__nand3_1 _28095_ (.A(_04114_),
    .B(_04112_),
    .C(_04110_),
    .Y(_04123_));
 sky130_fd_sc_hd__o21ai_2 _28096_ (.A1(_04113_),
    .A2(_04115_),
    .B1(net144),
    .Y(_04124_));
 sky130_fd_sc_hd__o211ai_1 _28097_ (.A1(net156),
    .A2(net154),
    .B1(_04122_),
    .C1(_04123_),
    .Y(_04125_));
 sky130_fd_sc_hd__o21ai_4 _28098_ (.A1(_04121_),
    .A2(_04124_),
    .B1(_04120_),
    .Y(_04126_));
 sky130_fd_sc_hd__o22a_4 _28099_ (.A1(net144),
    .A2(_04109_),
    .B1(_04121_),
    .B2(_04124_),
    .X(_04127_));
 sky130_fd_sc_hd__o211a_1 _28100_ (.A1(_04108_),
    .A2(net144),
    .B1(net197),
    .C1(_04119_),
    .X(_04129_));
 sky130_fd_sc_hd__o211ai_4 _28101_ (.A1(_04108_),
    .A2(net144),
    .B1(net197),
    .C1(_04119_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand3_2 _28102_ (.A(_04125_),
    .B(net201),
    .C(_04120_),
    .Y(_04131_));
 sky130_fd_sc_hd__and2_1 _28103_ (.A(_04130_),
    .B(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__nand2_1 _28104_ (.A(_04130_),
    .B(_04131_),
    .Y(_04133_));
 sky130_fd_sc_hd__nand4_1 _28105_ (.A(_03307_),
    .B(_03308_),
    .C(_03545_),
    .D(_03547_),
    .Y(_04134_));
 sky130_fd_sc_hd__a21oi_1 _28106_ (.A1(_07565_),
    .A2(_03762_),
    .B1(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__nor3_1 _28107_ (.A(_04134_),
    .B(_03771_),
    .C(_03769_),
    .Y(_04136_));
 sky130_fd_sc_hd__o211ai_2 _28108_ (.A1(_07565_),
    .A2(_03762_),
    .B1(_04135_),
    .C1(_03956_),
    .Y(_04137_));
 sky130_fd_sc_hd__o211ai_4 _28109_ (.A1(_03960_),
    .A2(_03955_),
    .B1(_03958_),
    .C1(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__nand4_4 _28110_ (.A(_04136_),
    .B(_03958_),
    .C(_03956_),
    .D(_03320_),
    .Y(_04140_));
 sky130_fd_sc_hd__nand2_2 _28111_ (.A(_04138_),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__a21oi_2 _28112_ (.A1(_04138_),
    .A2(_04140_),
    .B1(_04133_),
    .Y(_04142_));
 sky130_fd_sc_hd__a31o_1 _28113_ (.A1(_04133_),
    .A2(_04138_),
    .A3(_04140_),
    .B1(_09578_),
    .X(_04143_));
 sky130_fd_sc_hd__and3_1 _28114_ (.A(_04126_),
    .B(_09574_),
    .C(_09572_),
    .X(_04144_));
 sky130_fd_sc_hd__a22o_2 _28115_ (.A1(_04130_),
    .A2(_04131_),
    .B1(_04138_),
    .B2(_04140_),
    .X(_04145_));
 sky130_fd_sc_hd__o211ai_4 _28116_ (.A1(_04126_),
    .A2(net197),
    .B1(_04140_),
    .C1(_04138_),
    .Y(_04146_));
 sky130_fd_sc_hd__o2111ai_4 _28117_ (.A1(net197),
    .A2(_04126_),
    .B1(_04130_),
    .C1(_04138_),
    .D1(_04140_),
    .Y(_04147_));
 sky130_fd_sc_hd__o221ai_4 _28118_ (.A1(net142),
    .A2(_09573_),
    .B1(_04129_),
    .B2(_04146_),
    .C1(_04145_),
    .Y(_04148_));
 sky130_fd_sc_hd__a31o_2 _28119_ (.A1(net132),
    .A2(_04145_),
    .A3(_04147_),
    .B1(_04144_),
    .X(_04149_));
 sky130_fd_sc_hd__o22ai_4 _28120_ (.A1(net132),
    .A2(_04126_),
    .B1(_04142_),
    .B2(_04143_),
    .Y(_04151_));
 sky130_fd_sc_hd__a22oi_4 _28121_ (.A1(_03969_),
    .A2(_03951_),
    .B1(_03795_),
    .B2(_03783_),
    .Y(_04152_));
 sky130_fd_sc_hd__a21o_1 _28122_ (.A1(_03968_),
    .A2(_03971_),
    .B1(_03972_),
    .X(_04153_));
 sky130_fd_sc_hd__a21oi_2 _28123_ (.A1(_03968_),
    .A2(_03971_),
    .B1(_03972_),
    .Y(_04154_));
 sky130_fd_sc_hd__a311oi_4 _28124_ (.A1(net132),
    .A2(_04145_),
    .A3(_04147_),
    .B1(_04144_),
    .C1(_07936_),
    .Y(_04155_));
 sky130_fd_sc_hd__o211ai_4 _28125_ (.A1(net132),
    .A2(_04127_),
    .B1(_07935_),
    .C1(_04148_),
    .Y(_04156_));
 sky130_fd_sc_hd__o221ai_4 _28126_ (.A1(net132),
    .A2(_04126_),
    .B1(_04142_),
    .B2(_04143_),
    .C1(_07936_),
    .Y(_04157_));
 sky130_fd_sc_hd__nand2_1 _28127_ (.A(_04156_),
    .B(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__o211a_1 _28128_ (.A1(_03972_),
    .A2(_04152_),
    .B1(_04156_),
    .C1(_04157_),
    .X(_04159_));
 sky130_fd_sc_hd__o211ai_4 _28129_ (.A1(_03972_),
    .A2(_04152_),
    .B1(_04156_),
    .C1(_04157_),
    .Y(_04160_));
 sky130_fd_sc_hd__a21oi_1 _28130_ (.A1(_04156_),
    .A2(_04157_),
    .B1(_04153_),
    .Y(_04162_));
 sky130_fd_sc_hd__a21o_1 _28131_ (.A1(_04156_),
    .A2(_04157_),
    .B1(_04153_),
    .X(_04163_));
 sky130_fd_sc_hd__o22ai_2 _28132_ (.A1(net141),
    .A2(net139),
    .B1(_04159_),
    .B2(_04162_),
    .Y(_04164_));
 sky130_fd_sc_hd__or3_2 _28133_ (.A(net141),
    .B(net140),
    .C(_04151_),
    .X(_04165_));
 sky130_fd_sc_hd__inv_2 _28134_ (.A(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__o211ai_4 _28135_ (.A1(net141),
    .A2(net140),
    .B1(_04160_),
    .C1(_04163_),
    .Y(_04167_));
 sky130_fd_sc_hd__o31a_1 _28136_ (.A1(net141),
    .A2(net140),
    .A3(_04151_),
    .B1(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__inv_2 _28137_ (.A(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__a22oi_4 _28138_ (.A1(_07556_),
    .A2(_07558_),
    .B1(_04165_),
    .B2(_04167_),
    .Y(_04170_));
 sky130_fd_sc_hd__o221ai_4 _28139_ (.A1(net221),
    .A2(net219),
    .B1(net130),
    .B2(_04149_),
    .C1(_04164_),
    .Y(_04171_));
 sky130_fd_sc_hd__o21ai_1 _28140_ (.A1(_07560_),
    .A2(net217),
    .B1(_04167_),
    .Y(_04174_));
 sky130_fd_sc_hd__o311a_1 _28141_ (.A1(_10479_),
    .A2(_04159_),
    .A3(_04162_),
    .B1(_04165_),
    .C1(_07564_),
    .X(_04175_));
 sky130_fd_sc_hd__o211ai_4 _28142_ (.A1(net130),
    .A2(_04151_),
    .B1(_07564_),
    .C1(_04167_),
    .Y(_04176_));
 sky130_fd_sc_hd__o21a_1 _28143_ (.A1(_04166_),
    .A2(_04174_),
    .B1(_04171_),
    .X(_04177_));
 sky130_fd_sc_hd__o211ai_4 _28144_ (.A1(_06922_),
    .A2(_03799_),
    .B1(_03816_),
    .C1(_03990_),
    .Y(_04178_));
 sky130_fd_sc_hd__a32o_2 _28145_ (.A1(_03801_),
    .A2(_03816_),
    .A3(_03990_),
    .B1(_03985_),
    .B2(_03981_),
    .X(_04179_));
 sky130_fd_sc_hd__o211ai_2 _28146_ (.A1(_04174_),
    .A2(_04166_),
    .B1(_04171_),
    .C1(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__o221ai_4 _28147_ (.A1(net137),
    .A2(net135),
    .B1(_04179_),
    .B2(_04177_),
    .C1(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__or3_1 _28148_ (.A(net137),
    .B(net135),
    .C(_04168_),
    .X(_04182_));
 sky130_fd_sc_hd__o21ai_2 _28149_ (.A1(_04170_),
    .A2(_04175_),
    .B1(_04179_),
    .Y(_04183_));
 sky130_fd_sc_hd__a41oi_4 _28150_ (.A1(_03988_),
    .A2(_04171_),
    .A3(_04176_),
    .A4(_04178_),
    .B1(_10953_),
    .Y(_04185_));
 sky130_fd_sc_hd__nand2_1 _28151_ (.A(_04185_),
    .B(_04183_),
    .Y(_04186_));
 sky130_fd_sc_hd__o311a_1 _28152_ (.A1(net137),
    .A2(net135),
    .A3(_04168_),
    .B1(_11464_),
    .C1(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__a221oi_4 _28153_ (.A1(_10953_),
    .A2(_04169_),
    .B1(_04185_),
    .B2(_04183_),
    .C1(_07247_),
    .Y(_04188_));
 sky130_fd_sc_hd__o211ai_1 _28154_ (.A1(_10954_),
    .A2(_04168_),
    .B1(_07246_),
    .C1(_04186_),
    .Y(_04189_));
 sky130_fd_sc_hd__a2bb2oi_1 _28155_ (.A1_N(_07242_),
    .A2_N(net248),
    .B1(_04182_),
    .B2(_04186_),
    .Y(_04190_));
 sky130_fd_sc_hd__o211ai_4 _28156_ (.A1(_04169_),
    .A2(_10954_),
    .B1(_07247_),
    .C1(_04181_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand4_1 _28157_ (.A(_03999_),
    .B(_04013_),
    .C(_04189_),
    .D(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__o2bb2ai_1 _28158_ (.A1_N(_03999_),
    .A2_N(_04013_),
    .B1(_04188_),
    .B2(_04190_),
    .Y(_04193_));
 sky130_fd_sc_hd__o211a_1 _28159_ (.A1(_11459_),
    .A2(net129),
    .B1(_04192_),
    .C1(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__a31oi_1 _28160_ (.A1(_11465_),
    .A2(_04192_),
    .A3(_04193_),
    .B1(_04187_),
    .Y(_04196_));
 sky130_fd_sc_hd__and4_1 _28161_ (.A(_03382_),
    .B(_03383_),
    .C(_03617_),
    .D(_03618_),
    .X(_04197_));
 sky130_fd_sc_hd__nand4_1 _28162_ (.A(_04197_),
    .B(_04016_),
    .C(_03830_),
    .D(_03829_),
    .Y(_04198_));
 sky130_fd_sc_hd__o211ai_1 _28163_ (.A1(_04018_),
    .A2(_04015_),
    .B1(_04017_),
    .C1(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand4_1 _28164_ (.A(_04197_),
    .B(_03830_),
    .C(_03829_),
    .D(_03381_),
    .Y(_04200_));
 sky130_fd_sc_hd__nand3b_1 _28165_ (.A_N(_04200_),
    .B(_04017_),
    .C(_04016_),
    .Y(_04201_));
 sky130_fd_sc_hd__nand2_1 _28166_ (.A(_04199_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__o21ai_1 _28167_ (.A1(_04187_),
    .A2(_04194_),
    .B1(_06922_),
    .Y(_04203_));
 sky130_fd_sc_hd__and3_1 _28168_ (.A(_04196_),
    .B(_06921_),
    .C(_06919_),
    .X(_04204_));
 sky130_fd_sc_hd__o41a_1 _28169_ (.A1(_06918_),
    .A2(net249),
    .A3(_04187_),
    .A4(_04194_),
    .B1(_04203_),
    .X(_04205_));
 sky130_fd_sc_hd__inv_2 _28170_ (.A(_04205_),
    .Y(_04207_));
 sky130_fd_sc_hd__a21oi_1 _28171_ (.A1(_04202_),
    .A2(_04207_),
    .B1(_11944_),
    .Y(_04208_));
 sky130_fd_sc_hd__or2_1 _28172_ (.A(_04196_),
    .B(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__xnor2_1 _28173_ (.A(_04024_),
    .B(_04209_),
    .Y(net111));
 sky130_fd_sc_hd__o31ai_1 _28174_ (.A1(_03837_),
    .A2(_04021_),
    .A3(_04209_),
    .B1(_05119_),
    .Y(_04210_));
 sky130_fd_sc_hd__o311a_1 _28175_ (.A1(_03399_),
    .A2(net24),
    .A3(_10962_),
    .B1(_04030_),
    .C1(_04035_),
    .X(_04211_));
 sky130_fd_sc_hd__a31o_2 _28176_ (.A1(_11471_),
    .A2(_04030_),
    .A3(_04035_),
    .B1(_07550_),
    .X(_04212_));
 sky130_fd_sc_hd__a311oi_4 _28177_ (.A1(_11471_),
    .A2(_04030_),
    .A3(_04035_),
    .B1(_10970_),
    .C1(_07550_),
    .Y(_04213_));
 sky130_fd_sc_hd__o22a_1 _28178_ (.A1(_10965_),
    .A2(_10967_),
    .B1(_07550_),
    .B2(_04211_),
    .X(_04214_));
 sky130_fd_sc_hd__nor2_1 _28179_ (.A(_04213_),
    .B(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__o211ai_2 _28180_ (.A1(_03867_),
    .A2(net152),
    .B1(_04042_),
    .C1(_03881_),
    .Y(_04217_));
 sky130_fd_sc_hd__o221ai_4 _28181_ (.A1(_04213_),
    .A2(_04214_),
    .B1(_04043_),
    .B2(_04046_),
    .C1(_04042_),
    .Y(_04218_));
 sky130_fd_sc_hd__o211ai_4 _28182_ (.A1(_10492_),
    .A2(_04039_),
    .B1(_04215_),
    .C1(_04217_),
    .Y(_04219_));
 sky130_fd_sc_hd__o211ai_4 _28183_ (.A1(net183),
    .A2(net182),
    .B1(_04218_),
    .C1(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__and3_1 _28184_ (.A(_07913_),
    .B(_07915_),
    .C(_04212_),
    .X(_04221_));
 sky130_fd_sc_hd__a22oi_4 _28185_ (.A1(_07913_),
    .A2(_07915_),
    .B1(_04218_),
    .B2(_04219_),
    .Y(_04222_));
 sky130_fd_sc_hd__o21ai_4 _28186_ (.A1(_07916_),
    .A2(_04212_),
    .B1(_04220_),
    .Y(_04223_));
 sky130_fd_sc_hd__a211o_1 _28187_ (.A1(_07917_),
    .A2(_04212_),
    .B1(_04222_),
    .C1(net150),
    .X(_04224_));
 sky130_fd_sc_hd__o311a_1 _28188_ (.A1(_07550_),
    .A2(_07916_),
    .A3(_04211_),
    .B1(net150),
    .C1(_04220_),
    .X(_04225_));
 sky130_fd_sc_hd__o211ai_2 _28189_ (.A1(_07916_),
    .A2(_04212_),
    .B1(net150),
    .C1(_04220_),
    .Y(_04226_));
 sky130_fd_sc_hd__o41a_1 _28190_ (.A1(net164),
    .A2(_10490_),
    .A3(_04221_),
    .A4(_04222_),
    .B1(_04226_),
    .X(_04228_));
 sky130_fd_sc_hd__o41ai_4 _28191_ (.A1(net164),
    .A2(_10490_),
    .A3(_04221_),
    .A4(_04222_),
    .B1(_04226_),
    .Y(_04229_));
 sky130_fd_sc_hd__a21oi_1 _28192_ (.A1(_04066_),
    .A2(_04068_),
    .B1(_04057_),
    .Y(_04230_));
 sky130_fd_sc_hd__a31oi_4 _28193_ (.A1(_04060_),
    .A2(_04066_),
    .A3(_04068_),
    .B1(_04057_),
    .Y(_04231_));
 sky130_fd_sc_hd__o211a_1 _28194_ (.A1(net152),
    .A2(_04054_),
    .B1(_04072_),
    .C1(_04228_),
    .X(_04232_));
 sky130_fd_sc_hd__o21ai_2 _28195_ (.A1(_04228_),
    .A2(_04231_),
    .B1(net159),
    .Y(_04233_));
 sky130_fd_sc_hd__o211ai_2 _28196_ (.A1(net152),
    .A2(_04054_),
    .B1(_04072_),
    .C1(_04229_),
    .Y(_04234_));
 sky130_fd_sc_hd__or4_1 _28197_ (.A(net181),
    .B(net179),
    .C(_04221_),
    .D(_04222_),
    .X(_04235_));
 sky130_fd_sc_hd__o311ai_4 _28198_ (.A1(_04059_),
    .A2(_04229_),
    .A3(_04230_),
    .B1(_04234_),
    .C1(net159),
    .Y(_04236_));
 sky130_fd_sc_hd__o31a_2 _28199_ (.A1(net159),
    .A2(_04221_),
    .A3(_04222_),
    .B1(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__o221a_1 _28200_ (.A1(net159),
    .A2(_04223_),
    .B1(_04232_),
    .B2(_04233_),
    .C1(_10027_),
    .X(_04239_));
 sky130_fd_sc_hd__o221ai_4 _28201_ (.A1(net159),
    .A2(_04223_),
    .B1(_04232_),
    .B2(_04233_),
    .C1(_10027_),
    .Y(_04240_));
 sky130_fd_sc_hd__o211ai_4 _28202_ (.A1(net167),
    .A2(_10024_),
    .B1(_04235_),
    .C1(_04236_),
    .Y(_04241_));
 sky130_fd_sc_hd__nand2_1 _28203_ (.A(_04240_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__nand4_1 _28204_ (.A(_03485_),
    .B(_03486_),
    .C(_03712_),
    .D(_03714_),
    .Y(_04243_));
 sky130_fd_sc_hd__a211oi_2 _28205_ (.A1(_03890_),
    .A2(_03905_),
    .B1(_04243_),
    .C1(_03909_),
    .Y(_04244_));
 sky130_fd_sc_hd__nand2_1 _28206_ (.A(_04082_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__o211ai_4 _28207_ (.A1(_04087_),
    .A2(_04081_),
    .B1(_04083_),
    .C1(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__nand4_4 _28208_ (.A(_04244_),
    .B(_04083_),
    .C(_04082_),
    .D(_03495_),
    .Y(_04247_));
 sky130_fd_sc_hd__nand3_1 _28209_ (.A(_04242_),
    .B(_04246_),
    .C(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__a21o_1 _28210_ (.A1(_04246_),
    .A2(_04247_),
    .B1(_04242_),
    .X(_04250_));
 sky130_fd_sc_hd__a22o_1 _28211_ (.A1(_04240_),
    .A2(_04241_),
    .B1(_04246_),
    .B2(_04247_),
    .X(_04251_));
 sky130_fd_sc_hd__nand3_2 _28212_ (.A(_04241_),
    .B(_04246_),
    .C(_04247_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand4_2 _28213_ (.A(_04240_),
    .B(_04241_),
    .C(_04246_),
    .D(_04247_),
    .Y(_04253_));
 sky130_fd_sc_hd__nand3_2 _28214_ (.A(_04251_),
    .B(_04253_),
    .C(net149),
    .Y(_04254_));
 sky130_fd_sc_hd__o221a_1 _28215_ (.A1(net159),
    .A2(_04223_),
    .B1(_04232_),
    .B2(_04233_),
    .C1(_08715_),
    .X(_04255_));
 sky130_fd_sc_hd__or3_2 _28216_ (.A(net157),
    .B(_08712_),
    .C(_04237_),
    .X(_04256_));
 sky130_fd_sc_hd__o21ai_2 _28217_ (.A1(_08705_),
    .A2(_08707_),
    .B1(_04237_),
    .Y(_04257_));
 sky130_fd_sc_hd__nand3_1 _28218_ (.A(_04250_),
    .B(net149),
    .C(_04248_),
    .Y(_04258_));
 sky130_fd_sc_hd__a31o_2 _28219_ (.A1(_04251_),
    .A2(_04253_),
    .A3(net149),
    .B1(_04255_),
    .X(_04259_));
 sky130_fd_sc_hd__and3_1 _28220_ (.A(_04258_),
    .B(_09124_),
    .C(_04257_),
    .X(_04261_));
 sky130_fd_sc_hd__a211o_2 _28221_ (.A1(_04254_),
    .A2(_04256_),
    .B1(net148),
    .C1(net147),
    .X(_04262_));
 sky130_fd_sc_hd__a311oi_2 _28222_ (.A1(_04251_),
    .A2(_04253_),
    .A3(net149),
    .B1(_04255_),
    .C1(net171),
    .Y(_04263_));
 sky130_fd_sc_hd__nand3_4 _28223_ (.A(_04254_),
    .B(_04256_),
    .C(_09594_),
    .Y(_04264_));
 sky130_fd_sc_hd__o211ai_4 _28224_ (.A1(net189),
    .A2(net186),
    .B1(_04257_),
    .C1(_04258_),
    .Y(_04265_));
 sky130_fd_sc_hd__o221a_1 _28225_ (.A1(_03922_),
    .A2(_03923_),
    .B1(_04091_),
    .B2(_09139_),
    .C1(_03920_),
    .X(_04266_));
 sky130_fd_sc_hd__a31o_1 _28226_ (.A1(_03921_),
    .A2(_04094_),
    .A3(_04098_),
    .B1(_04099_),
    .X(_04267_));
 sky130_fd_sc_hd__a31oi_2 _28227_ (.A1(_03921_),
    .A2(_04094_),
    .A3(_04098_),
    .B1(_04099_),
    .Y(_04268_));
 sky130_fd_sc_hd__a21oi_1 _28228_ (.A1(_04264_),
    .A2(_04265_),
    .B1(_04267_),
    .Y(_04269_));
 sky130_fd_sc_hd__o2bb2ai_4 _28229_ (.A1_N(_04264_),
    .A2_N(_04265_),
    .B1(_04266_),
    .B2(_04097_),
    .Y(_04270_));
 sky130_fd_sc_hd__and3_1 _28230_ (.A(_04264_),
    .B(_04265_),
    .C(_04267_),
    .X(_04272_));
 sky130_fd_sc_hd__nand3_1 _28231_ (.A(_04264_),
    .B(_04265_),
    .C(_04267_),
    .Y(_04273_));
 sky130_fd_sc_hd__a31oi_4 _28232_ (.A1(_04264_),
    .A2(_04265_),
    .A3(_04267_),
    .B1(_09124_),
    .Y(_04274_));
 sky130_fd_sc_hd__nand3_2 _28233_ (.A(net145),
    .B(_04270_),
    .C(_04273_),
    .Y(_04275_));
 sky130_fd_sc_hd__o22ai_2 _28234_ (.A1(net148),
    .A2(net147),
    .B1(_04269_),
    .B2(_04272_),
    .Y(_04276_));
 sky130_fd_sc_hd__a21oi_2 _28235_ (.A1(_04274_),
    .A2(_04270_),
    .B1(_04261_),
    .Y(_04277_));
 sky130_fd_sc_hd__a311o_1 _28236_ (.A1(net145),
    .A2(_04270_),
    .A3(_04273_),
    .B1(net144),
    .C1(_04261_),
    .X(_04278_));
 sky130_fd_sc_hd__o221ai_4 _28237_ (.A1(net201),
    .A2(_03927_),
    .B1(net178),
    .B2(_04109_),
    .C1(_03946_),
    .Y(_04279_));
 sky130_fd_sc_hd__a31oi_2 _28238_ (.A1(_03933_),
    .A2(_03946_),
    .A3(_04110_),
    .B1(_04111_),
    .Y(_04280_));
 sky130_fd_sc_hd__a21oi_1 _28239_ (.A1(_04274_),
    .A2(_04270_),
    .B1(_09140_),
    .Y(_04281_));
 sky130_fd_sc_hd__a221oi_4 _28240_ (.A1(_09124_),
    .A2(_04259_),
    .B1(_04274_),
    .B2(_04270_),
    .C1(_09140_),
    .Y(_04284_));
 sky130_fd_sc_hd__nand3_2 _28241_ (.A(_04275_),
    .B(_09139_),
    .C(_04262_),
    .Y(_04285_));
 sky130_fd_sc_hd__a2bb2oi_4 _28242_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_04262_),
    .B2(_04275_),
    .Y(_04286_));
 sky130_fd_sc_hd__o221ai_4 _28243_ (.A1(net194),
    .A2(net190),
    .B1(_04259_),
    .B2(net145),
    .C1(_04276_),
    .Y(_04287_));
 sky130_fd_sc_hd__o2111ai_1 _28244_ (.A1(_04113_),
    .A2(_04115_),
    .B1(_04285_),
    .C1(_04287_),
    .D1(_04110_),
    .Y(_04288_));
 sky130_fd_sc_hd__o21ai_1 _28245_ (.A1(_04284_),
    .A2(_04286_),
    .B1(_04280_),
    .Y(_04289_));
 sky130_fd_sc_hd__o211ai_2 _28246_ (.A1(net156),
    .A2(net154),
    .B1(_04288_),
    .C1(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__a211o_1 _28247_ (.A1(_04262_),
    .A2(_04275_),
    .B1(net156),
    .C1(net154),
    .X(_04291_));
 sky130_fd_sc_hd__inv_2 _28248_ (.A(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__nand3_2 _28249_ (.A(_04280_),
    .B(_04285_),
    .C(_04287_),
    .Y(_04293_));
 sky130_fd_sc_hd__o2bb2ai_2 _28250_ (.A1_N(_04112_),
    .A2_N(_04279_),
    .B1(_04284_),
    .B2(_04286_),
    .Y(_04295_));
 sky130_fd_sc_hd__o211ai_2 _28251_ (.A1(net156),
    .A2(net154),
    .B1(_04293_),
    .C1(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hd__a31o_2 _28252_ (.A1(net144),
    .A2(_04293_),
    .A3(_04295_),
    .B1(_04292_),
    .X(_04297_));
 sky130_fd_sc_hd__a31oi_4 _28253_ (.A1(net144),
    .A2(_04293_),
    .A3(_04295_),
    .B1(_04292_),
    .Y(_04298_));
 sky130_fd_sc_hd__o211ai_4 _28254_ (.A1(_08724_),
    .A2(net196),
    .B1(_04278_),
    .C1(_04290_),
    .Y(_04299_));
 sky130_fd_sc_hd__o211ai_4 _28255_ (.A1(net144),
    .A2(_04277_),
    .B1(net178),
    .C1(_04296_),
    .Y(_04300_));
 sky130_fd_sc_hd__and2_1 _28256_ (.A(_04299_),
    .B(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__nand2_2 _28257_ (.A(_04299_),
    .B(_04300_),
    .Y(_04302_));
 sky130_fd_sc_hd__o2bb2ai_2 _28258_ (.A1_N(_04138_),
    .A2_N(_04140_),
    .B1(net201),
    .B2(_04127_),
    .Y(_04303_));
 sky130_fd_sc_hd__a31oi_2 _28259_ (.A1(_04131_),
    .A2(_04138_),
    .A3(_04140_),
    .B1(_04129_),
    .Y(_04304_));
 sky130_fd_sc_hd__o311a_2 _28260_ (.A1(_08311_),
    .A2(net215),
    .A3(_04127_),
    .B1(_04146_),
    .C1(_04302_),
    .X(_04306_));
 sky130_fd_sc_hd__o211ai_2 _28261_ (.A1(net201),
    .A2(_04127_),
    .B1(_04146_),
    .C1(_04302_),
    .Y(_04307_));
 sky130_fd_sc_hd__o2111ai_4 _28262_ (.A1(net197),
    .A2(_04126_),
    .B1(_04299_),
    .C1(_04300_),
    .D1(_04303_),
    .Y(_04308_));
 sky130_fd_sc_hd__o22ai_4 _28263_ (.A1(net142),
    .A2(_09573_),
    .B1(_04302_),
    .B2(_04304_),
    .Y(_04309_));
 sky130_fd_sc_hd__o211ai_4 _28264_ (.A1(net142),
    .A2(_09573_),
    .B1(_04307_),
    .C1(_04308_),
    .Y(_04310_));
 sky130_fd_sc_hd__or3_2 _28265_ (.A(net142),
    .B(_09573_),
    .C(_04298_),
    .X(_04311_));
 sky130_fd_sc_hd__o32a_1 _28266_ (.A1(net142),
    .A2(_09573_),
    .A3(_04298_),
    .B1(_04306_),
    .B2(_04309_),
    .X(_04312_));
 sky130_fd_sc_hd__o22ai_4 _28267_ (.A1(net132),
    .A2(_04298_),
    .B1(_04306_),
    .B2(_04309_),
    .Y(_04313_));
 sky130_fd_sc_hd__a21oi_4 _28268_ (.A1(_04310_),
    .A2(_04311_),
    .B1(net201),
    .Y(_04314_));
 sky130_fd_sc_hd__a22o_2 _28269_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_04310_),
    .B2(_04311_),
    .X(_04315_));
 sky130_fd_sc_hd__o22a_1 _28270_ (.A1(_08311_),
    .A2(net215),
    .B1(_04306_),
    .B2(_04309_),
    .X(_04317_));
 sky130_fd_sc_hd__o221a_1 _28271_ (.A1(net132),
    .A2(_04298_),
    .B1(_04306_),
    .B2(_04309_),
    .C1(net201),
    .X(_04318_));
 sky130_fd_sc_hd__o221ai_4 _28272_ (.A1(_08311_),
    .A2(net215),
    .B1(net132),
    .B2(_04298_),
    .C1(_04310_),
    .Y(_04319_));
 sky130_fd_sc_hd__a21oi_1 _28273_ (.A1(_04311_),
    .A2(_04317_),
    .B1(_04314_),
    .Y(_04320_));
 sky130_fd_sc_hd__nand2_1 _28274_ (.A(_04315_),
    .B(_04319_),
    .Y(_04321_));
 sky130_fd_sc_hd__and4_1 _28275_ (.A(_03560_),
    .B(_03563_),
    .C(_03783_),
    .D(_03785_),
    .X(_04322_));
 sky130_fd_sc_hd__nand4_2 _28276_ (.A(_03560_),
    .B(_03563_),
    .C(_03783_),
    .D(_03785_),
    .Y(_04323_));
 sky130_fd_sc_hd__a211oi_4 _28277_ (.A1(_03951_),
    .A2(_03969_),
    .B1(_04323_),
    .C1(_03972_),
    .Y(_04324_));
 sky130_fd_sc_hd__nand3_1 _28278_ (.A(_04156_),
    .B(_04322_),
    .C(_03974_),
    .Y(_04325_));
 sky130_fd_sc_hd__a32oi_4 _28279_ (.A1(_04149_),
    .A2(_07934_),
    .A3(_07933_),
    .B1(_04324_),
    .B2(_04156_),
    .Y(_04326_));
 sky130_fd_sc_hd__o211a_1 _28280_ (.A1(_04154_),
    .A2(_04155_),
    .B1(_04157_),
    .C1(_04325_),
    .X(_04328_));
 sky130_fd_sc_hd__o211ai_4 _28281_ (.A1(_04154_),
    .A2(_04155_),
    .B1(_04157_),
    .C1(_04325_),
    .Y(_04329_));
 sky130_fd_sc_hd__nand4_2 _28282_ (.A(_04322_),
    .B(_03973_),
    .C(_03971_),
    .D(_03575_),
    .Y(_04330_));
 sky130_fd_sc_hd__nand4_4 _28283_ (.A(_04324_),
    .B(_04157_),
    .C(_04156_),
    .D(_03575_),
    .Y(_04331_));
 sky130_fd_sc_hd__a41o_1 _28284_ (.A1(_03575_),
    .A2(_04156_),
    .A3(_04157_),
    .A4(_04324_),
    .B1(_04328_),
    .X(_04332_));
 sky130_fd_sc_hd__a21oi_2 _28285_ (.A1(_04329_),
    .A2(_04331_),
    .B1(_04321_),
    .Y(_04333_));
 sky130_fd_sc_hd__o221ai_2 _28286_ (.A1(_04158_),
    .A2(_04330_),
    .B1(_04318_),
    .B2(_04314_),
    .C1(_04329_),
    .Y(_04334_));
 sky130_fd_sc_hd__o21ai_2 _28287_ (.A1(net141),
    .A2(net139),
    .B1(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__or3_2 _28288_ (.A(net141),
    .B(net139),
    .C(_04312_),
    .X(_04336_));
 sky130_fd_sc_hd__a22oi_1 _28289_ (.A1(_04315_),
    .A2(_04319_),
    .B1(_04329_),
    .B2(_04331_),
    .Y(_04337_));
 sky130_fd_sc_hd__a22o_1 _28290_ (.A1(_04315_),
    .A2(_04319_),
    .B1(_04329_),
    .B2(_04331_),
    .X(_04339_));
 sky130_fd_sc_hd__o22ai_4 _28291_ (.A1(net197),
    .A2(_04313_),
    .B1(_04330_),
    .B2(_04158_),
    .Y(_04340_));
 sky130_fd_sc_hd__a21oi_2 _28292_ (.A1(_04160_),
    .A2(_04326_),
    .B1(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__nand3_2 _28293_ (.A(_04319_),
    .B(_04329_),
    .C(_04331_),
    .Y(_04342_));
 sky130_fd_sc_hd__a211oi_1 _28294_ (.A1(_04326_),
    .A2(_04160_),
    .B1(_04314_),
    .C1(_04340_),
    .Y(_04343_));
 sky130_fd_sc_hd__o221ai_4 _28295_ (.A1(net141),
    .A2(net139),
    .B1(_04314_),
    .B2(_04342_),
    .C1(_04339_),
    .Y(_04344_));
 sky130_fd_sc_hd__o22a_1 _28296_ (.A1(net130),
    .A2(_04313_),
    .B1(_04333_),
    .B2(_04335_),
    .X(_04345_));
 sky130_fd_sc_hd__o211a_1 _28297_ (.A1(_03983_),
    .A2(_07247_),
    .B1(_04178_),
    .C1(_04176_),
    .X(_04346_));
 sky130_fd_sc_hd__a31o_1 _28298_ (.A1(_03988_),
    .A2(_04176_),
    .A3(_04178_),
    .B1(_04170_),
    .X(_04347_));
 sky130_fd_sc_hd__a31oi_2 _28299_ (.A1(_03988_),
    .A2(_04176_),
    .A3(_04178_),
    .B1(_04170_),
    .Y(_04348_));
 sky130_fd_sc_hd__o311a_1 _28300_ (.A1(_10479_),
    .A2(_04337_),
    .A3(_04343_),
    .B1(_04336_),
    .C1(_07935_),
    .X(_04350_));
 sky130_fd_sc_hd__nand3_4 _28301_ (.A(_04344_),
    .B(_07935_),
    .C(_04336_),
    .Y(_04351_));
 sky130_fd_sc_hd__o221a_1 _28302_ (.A1(net130),
    .A2(_04313_),
    .B1(_04333_),
    .B2(_04335_),
    .C1(_07936_),
    .X(_04352_));
 sky130_fd_sc_hd__o221ai_4 _28303_ (.A1(net130),
    .A2(_04313_),
    .B1(_04333_),
    .B2(_04335_),
    .C1(_07936_),
    .Y(_04353_));
 sky130_fd_sc_hd__o211a_1 _28304_ (.A1(_04170_),
    .A2(_04346_),
    .B1(_04351_),
    .C1(_04353_),
    .X(_04354_));
 sky130_fd_sc_hd__o211ai_2 _28305_ (.A1(_04170_),
    .A2(_04346_),
    .B1(_04351_),
    .C1(_04353_),
    .Y(_04355_));
 sky130_fd_sc_hd__a21oi_1 _28306_ (.A1(_04351_),
    .A2(_04353_),
    .B1(_04347_),
    .Y(_04356_));
 sky130_fd_sc_hd__a21o_1 _28307_ (.A1(_04351_),
    .A2(_04353_),
    .B1(_04347_),
    .X(_04357_));
 sky130_fd_sc_hd__o22ai_2 _28308_ (.A1(net137),
    .A2(net134),
    .B1(_04354_),
    .B2(_04356_),
    .Y(_04358_));
 sky130_fd_sc_hd__a211o_1 _28309_ (.A1(_04336_),
    .A2(_04344_),
    .B1(net137),
    .C1(net134),
    .X(_04359_));
 sky130_fd_sc_hd__o211ai_2 _28310_ (.A1(net137),
    .A2(net134),
    .B1(_04355_),
    .C1(_04357_),
    .Y(_04361_));
 sky130_fd_sc_hd__nand2_1 _28311_ (.A(_04359_),
    .B(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__o221a_1 _28312_ (.A1(net221),
    .A2(net219),
    .B1(_10954_),
    .B2(_04345_),
    .C1(_04358_),
    .X(_04363_));
 sky130_fd_sc_hd__o221ai_4 _28313_ (.A1(net221),
    .A2(net219),
    .B1(_10954_),
    .B2(_04345_),
    .C1(_04358_),
    .Y(_04364_));
 sky130_fd_sc_hd__o211ai_4 _28314_ (.A1(_07560_),
    .A2(net217),
    .B1(_04359_),
    .C1(_04361_),
    .Y(_04365_));
 sky130_fd_sc_hd__inv_2 _28315_ (.A(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__a31oi_4 _28316_ (.A1(_03999_),
    .A2(_04013_),
    .A3(_04191_),
    .B1(_04188_),
    .Y(_04367_));
 sky130_fd_sc_hd__a21o_1 _28317_ (.A1(_04364_),
    .A2(_04365_),
    .B1(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__a31oi_2 _28318_ (.A1(_04367_),
    .A2(_04365_),
    .A3(_04364_),
    .B1(_11464_),
    .Y(_04369_));
 sky130_fd_sc_hd__a32o_1 _28319_ (.A1(_11460_),
    .A2(_11462_),
    .A3(_04362_),
    .B1(_04369_),
    .B2(_04368_),
    .X(_04370_));
 sky130_fd_sc_hd__o21ai_1 _28320_ (.A1(_07242_),
    .A2(net248),
    .B1(_04370_),
    .Y(_04372_));
 sky130_fd_sc_hd__a221oi_1 _28321_ (.A1(_11464_),
    .A2(_04362_),
    .B1(_04369_),
    .B2(_04368_),
    .C1(_07247_),
    .Y(_04373_));
 sky130_fd_sc_hd__a221o_1 _28322_ (.A1(_11464_),
    .A2(_04362_),
    .B1(_04369_),
    .B2(_04368_),
    .C1(_07247_),
    .X(_04374_));
 sky130_fd_sc_hd__a31oi_1 _28323_ (.A1(_04199_),
    .A2(_04201_),
    .A3(_04203_),
    .B1(_04204_),
    .Y(_04375_));
 sky130_fd_sc_hd__a21boi_1 _28324_ (.A1(_04372_),
    .A2(_04374_),
    .B1_N(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__o21ba_1 _28325_ (.A1(_11944_),
    .A2(_04376_),
    .B1_N(_04370_),
    .X(_04377_));
 sky130_fd_sc_hd__xor2_1 _28326_ (.A(_04210_),
    .B(_04377_),
    .X(net112));
 sky130_fd_sc_hd__nor4b_1 _28327_ (.A(_03837_),
    .B(_04021_),
    .C(_04209_),
    .D_N(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__o211ai_2 _28328_ (.A1(_04212_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_04219_),
    .Y(_04379_));
 sky130_fd_sc_hd__o21ai_1 _28329_ (.A1(net183),
    .A2(net182),
    .B1(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__and3_2 _28330_ (.A(_04379_),
    .B(_07916_),
    .C(_08301_),
    .X(_04382_));
 sky130_fd_sc_hd__inv_2 _28331_ (.A(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__and3_1 _28332_ (.A(_04379_),
    .B(_07916_),
    .C(_10971_),
    .X(_04384_));
 sky130_fd_sc_hd__o2bb2a_1 _28333_ (.A1_N(_07916_),
    .A2_N(_04379_),
    .B1(_10967_),
    .B2(_10965_),
    .X(_04385_));
 sky130_fd_sc_hd__nor2_1 _28334_ (.A(_04384_),
    .B(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__o211ai_2 _28335_ (.A1(net152),
    .A2(_04054_),
    .B1(_04072_),
    .C1(_04224_),
    .Y(_04387_));
 sky130_fd_sc_hd__o221ai_4 _28336_ (.A1(_04384_),
    .A2(_04385_),
    .B1(_04225_),
    .B2(_04231_),
    .C1(_04224_),
    .Y(_04388_));
 sky130_fd_sc_hd__o211ai_4 _28337_ (.A1(_10492_),
    .A2(_04223_),
    .B1(_04386_),
    .C1(_04387_),
    .Y(_04389_));
 sky130_fd_sc_hd__o211ai_1 _28338_ (.A1(net181),
    .A2(net179),
    .B1(_04388_),
    .C1(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__a31o_4 _28339_ (.A1(_04388_),
    .A2(_04389_),
    .A3(net159),
    .B1(_04382_),
    .X(_04391_));
 sky130_fd_sc_hd__a21oi_1 _28340_ (.A1(_04383_),
    .A2(_04390_),
    .B1(_10491_),
    .Y(_04394_));
 sky130_fd_sc_hd__a2bb2o_2 _28341_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_04383_),
    .B2(_04390_),
    .X(_04395_));
 sky130_fd_sc_hd__a31o_1 _28342_ (.A1(_04388_),
    .A2(_04389_),
    .A3(net159),
    .B1(_10492_),
    .X(_04396_));
 sky130_fd_sc_hd__and3_2 _28343_ (.A(_04390_),
    .B(_10491_),
    .C(_04383_),
    .X(_04397_));
 sky130_fd_sc_hd__o2bb2ai_1 _28344_ (.A1_N(_04246_),
    .A2_N(_04247_),
    .B1(net152),
    .B2(_04237_),
    .Y(_04398_));
 sky130_fd_sc_hd__a31oi_2 _28345_ (.A1(_04241_),
    .A2(_04246_),
    .A3(_04247_),
    .B1(_04239_),
    .Y(_04399_));
 sky130_fd_sc_hd__o2111ai_4 _28346_ (.A1(_04382_),
    .A2(_04396_),
    .B1(_04395_),
    .C1(_04240_),
    .D1(_04252_),
    .Y(_04400_));
 sky130_fd_sc_hd__o211ai_2 _28347_ (.A1(_04394_),
    .A2(_04397_),
    .B1(_04398_),
    .C1(_04241_),
    .Y(_04401_));
 sky130_fd_sc_hd__o2111ai_2 _28348_ (.A1(_04396_),
    .A2(_04382_),
    .B1(_04241_),
    .C1(_04395_),
    .D1(_04398_),
    .Y(_04402_));
 sky130_fd_sc_hd__o211ai_2 _28349_ (.A1(_04394_),
    .A2(_04397_),
    .B1(_04240_),
    .C1(_04252_),
    .Y(_04403_));
 sky130_fd_sc_hd__o211ai_4 _28350_ (.A1(net157),
    .A2(_08712_),
    .B1(_04400_),
    .C1(_04401_),
    .Y(_04405_));
 sky130_fd_sc_hd__and3_1 _28351_ (.A(_08710_),
    .B(_08713_),
    .C(_04391_),
    .X(_04406_));
 sky130_fd_sc_hd__nand3_1 _28352_ (.A(_04402_),
    .B(_04403_),
    .C(net149),
    .Y(_04407_));
 sky130_fd_sc_hd__a31o_2 _28353_ (.A1(_04402_),
    .A2(_04403_),
    .A3(net149),
    .B1(_04406_),
    .X(_04408_));
 sky130_fd_sc_hd__o21ai_4 _28354_ (.A1(net149),
    .A2(_04391_),
    .B1(_04405_),
    .Y(_04409_));
 sky130_fd_sc_hd__o311a_1 _28355_ (.A1(net157),
    .A2(_08712_),
    .A3(_04391_),
    .B1(_09124_),
    .C1(_04405_),
    .X(_04410_));
 sky130_fd_sc_hd__o311a_1 _28356_ (.A1(net157),
    .A2(_04391_),
    .A3(_08712_),
    .B1(_10027_),
    .C1(_04405_),
    .X(_04411_));
 sky130_fd_sc_hd__o211ai_4 _28357_ (.A1(_04391_),
    .A2(net149),
    .B1(_10027_),
    .C1(_04405_),
    .Y(_04412_));
 sky130_fd_sc_hd__nand3b_1 _28358_ (.A_N(_04406_),
    .B(_04407_),
    .C(net152),
    .Y(_04413_));
 sky130_fd_sc_hd__nand2_1 _28359_ (.A(_04412_),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__nand4_1 _28360_ (.A(_03726_),
    .B(_03727_),
    .C(_03920_),
    .D(_03921_),
    .Y(_04416_));
 sky130_fd_sc_hd__a211oi_2 _28361_ (.A1(_04080_),
    .A2(_04096_),
    .B1(_04416_),
    .C1(_04099_),
    .Y(_04417_));
 sky130_fd_sc_hd__nand2_1 _28362_ (.A(_04264_),
    .B(_04417_),
    .Y(_04418_));
 sky130_fd_sc_hd__o211ai_4 _28363_ (.A1(_04268_),
    .A2(_04263_),
    .B1(_04265_),
    .C1(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__nand4_4 _28364_ (.A(_04417_),
    .B(_04265_),
    .C(_04264_),
    .D(_03736_),
    .Y(_04420_));
 sky130_fd_sc_hd__nand3_1 _28365_ (.A(_04414_),
    .B(_04419_),
    .C(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__a21o_1 _28366_ (.A1(_04419_),
    .A2(_04420_),
    .B1(_04414_),
    .X(_04422_));
 sky130_fd_sc_hd__a22o_1 _28367_ (.A1(_04412_),
    .A2(_04413_),
    .B1(_04419_),
    .B2(_04420_),
    .X(_04423_));
 sky130_fd_sc_hd__o211ai_4 _28368_ (.A1(_04408_),
    .A2(_10027_),
    .B1(_04420_),
    .C1(_04419_),
    .Y(_04424_));
 sky130_fd_sc_hd__nand4_1 _28369_ (.A(_04412_),
    .B(_04413_),
    .C(_04419_),
    .D(_04420_),
    .Y(_04425_));
 sky130_fd_sc_hd__o221ai_4 _28370_ (.A1(net148),
    .A2(net147),
    .B1(_04411_),
    .B2(_04424_),
    .C1(_04423_),
    .Y(_04427_));
 sky130_fd_sc_hd__a311o_1 _28371_ (.A1(_04402_),
    .A2(_04403_),
    .A3(net149),
    .B1(_04406_),
    .C1(net145),
    .X(_04428_));
 sky130_fd_sc_hd__o211ai_4 _28372_ (.A1(net148),
    .A2(net147),
    .B1(_04421_),
    .C1(_04422_),
    .Y(_04429_));
 sky130_fd_sc_hd__a31o_1 _28373_ (.A1(net145),
    .A2(_04423_),
    .A3(_04425_),
    .B1(_04410_),
    .X(_04430_));
 sky130_fd_sc_hd__and3_2 _28374_ (.A(_04429_),
    .B(_09562_),
    .C(_04428_),
    .X(_04431_));
 sky130_fd_sc_hd__o21ai_2 _28375_ (.A1(_09559_),
    .A2(_09560_),
    .B1(_04430_),
    .Y(_04432_));
 sky130_fd_sc_hd__a311oi_2 _28376_ (.A1(net145),
    .A2(_04423_),
    .A3(_04425_),
    .B1(net171),
    .C1(_04410_),
    .Y(_04433_));
 sky130_fd_sc_hd__o211ai_4 _28377_ (.A1(net145),
    .A2(_04409_),
    .B1(_09594_),
    .C1(_04427_),
    .Y(_04434_));
 sky130_fd_sc_hd__o211ai_4 _28378_ (.A1(_04408_),
    .A2(net145),
    .B1(net171),
    .C1(_04429_),
    .Y(_04435_));
 sky130_fd_sc_hd__o221a_1 _28379_ (.A1(_04111_),
    .A2(_04115_),
    .B1(_04277_),
    .B2(_09139_),
    .C1(_04110_),
    .X(_04436_));
 sky130_fd_sc_hd__o211a_1 _28380_ (.A1(_04108_),
    .A2(net176),
    .B1(_04285_),
    .C1(_04279_),
    .X(_04438_));
 sky130_fd_sc_hd__a31o_1 _28381_ (.A1(_04112_),
    .A2(_04279_),
    .A3(_04285_),
    .B1(_04286_),
    .X(_04439_));
 sky130_fd_sc_hd__a21oi_2 _28382_ (.A1(_04280_),
    .A2(_04285_),
    .B1(_04286_),
    .Y(_04440_));
 sky130_fd_sc_hd__a21oi_1 _28383_ (.A1(_04434_),
    .A2(_04435_),
    .B1(_04439_),
    .Y(_04441_));
 sky130_fd_sc_hd__o2bb2ai_4 _28384_ (.A1_N(_04434_),
    .A2_N(_04435_),
    .B1(_04436_),
    .B2(_04284_),
    .Y(_04442_));
 sky130_fd_sc_hd__o211a_1 _28385_ (.A1(_04286_),
    .A2(_04438_),
    .B1(_04435_),
    .C1(_04434_),
    .X(_04443_));
 sky130_fd_sc_hd__o211ai_4 _28386_ (.A1(_04286_),
    .A2(_04438_),
    .B1(_04435_),
    .C1(_04434_),
    .Y(_04444_));
 sky130_fd_sc_hd__nand3_1 _28387_ (.A(net144),
    .B(_04442_),
    .C(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__o22ai_2 _28388_ (.A1(net156),
    .A2(net154),
    .B1(_04441_),
    .B2(_04443_),
    .Y(_04446_));
 sky130_fd_sc_hd__a31oi_4 _28389_ (.A1(net144),
    .A2(_04442_),
    .A3(_04444_),
    .B1(_04431_),
    .Y(_04447_));
 sky130_fd_sc_hd__a31o_1 _28390_ (.A1(net144),
    .A2(_04442_),
    .A3(_04444_),
    .B1(_04431_),
    .X(_04449_));
 sky130_fd_sc_hd__o221ai_4 _28391_ (.A1(net201),
    .A2(_04127_),
    .B1(net178),
    .B2(_04298_),
    .C1(_04146_),
    .Y(_04450_));
 sky130_fd_sc_hd__o221ai_2 _28392_ (.A1(net197),
    .A2(_04126_),
    .B1(_04297_),
    .B2(net176),
    .C1(_04303_),
    .Y(_04451_));
 sky130_fd_sc_hd__a31oi_1 _28393_ (.A1(net144),
    .A2(_04442_),
    .A3(_04444_),
    .B1(_09140_),
    .Y(_04452_));
 sky130_fd_sc_hd__a311oi_4 _28394_ (.A1(net144),
    .A2(_04442_),
    .A3(_04444_),
    .B1(_04431_),
    .C1(_09140_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand3_2 _28395_ (.A(_04445_),
    .B(_09139_),
    .C(_04432_),
    .Y(_04454_));
 sky130_fd_sc_hd__a2bb2oi_2 _28396_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_04432_),
    .B2(_04445_),
    .Y(_04455_));
 sky130_fd_sc_hd__o221ai_4 _28397_ (.A1(net194),
    .A2(net190),
    .B1(net144),
    .B2(_04430_),
    .C1(_04446_),
    .Y(_04456_));
 sky130_fd_sc_hd__o2111ai_1 _28398_ (.A1(_04298_),
    .A2(net178),
    .B1(_04454_),
    .C1(_04451_),
    .D1(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__o2bb2ai_1 _28399_ (.A1_N(_04299_),
    .A2_N(_04451_),
    .B1(_04453_),
    .B2(_04455_),
    .Y(_04458_));
 sky130_fd_sc_hd__o211ai_2 _28400_ (.A1(net142),
    .A2(_09573_),
    .B1(_04457_),
    .C1(_04458_),
    .Y(_04460_));
 sky130_fd_sc_hd__o221ai_4 _28401_ (.A1(_04297_),
    .A2(net176),
    .B1(_09139_),
    .B2(_04447_),
    .C1(_04450_),
    .Y(_04461_));
 sky130_fd_sc_hd__o2bb2ai_1 _28402_ (.A1_N(_04300_),
    .A2_N(_04450_),
    .B1(_04453_),
    .B2(_04455_),
    .Y(_04462_));
 sky130_fd_sc_hd__o221ai_4 _28403_ (.A1(net142),
    .A2(_09573_),
    .B1(_04453_),
    .B2(_04461_),
    .C1(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__o21ai_4 _28404_ (.A1(net132),
    .A2(_04447_),
    .B1(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__inv_2 _28405_ (.A(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__o211ai_4 _28406_ (.A1(net132),
    .A2(_04449_),
    .B1(_04460_),
    .C1(net176),
    .Y(_04466_));
 sky130_fd_sc_hd__o211a_1 _28407_ (.A1(net132),
    .A2(_04447_),
    .B1(net178),
    .C1(_04463_),
    .X(_04467_));
 sky130_fd_sc_hd__o211ai_2 _28408_ (.A1(net132),
    .A2(_04447_),
    .B1(net178),
    .C1(_04463_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand2_2 _28409_ (.A(_04466_),
    .B(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hd__a31oi_4 _28410_ (.A1(_04319_),
    .A2(_04329_),
    .A3(_04331_),
    .B1(_04314_),
    .Y(_04471_));
 sky130_fd_sc_hd__o21ai_1 _28411_ (.A1(_04314_),
    .A2(_04341_),
    .B1(_04469_),
    .Y(_04472_));
 sky130_fd_sc_hd__o311ai_4 _28412_ (.A1(_04314_),
    .A2(_04469_),
    .A3(_04341_),
    .B1(net130),
    .C1(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__o311a_2 _28413_ (.A1(_08311_),
    .A2(net215),
    .A3(_04312_),
    .B1(_04342_),
    .C1(_04469_),
    .X(_04474_));
 sky130_fd_sc_hd__o22ai_4 _28414_ (.A1(net141),
    .A2(net139),
    .B1(_04469_),
    .B2(_04471_),
    .Y(_04475_));
 sky130_fd_sc_hd__o22ai_4 _28415_ (.A1(net130),
    .A2(_04465_),
    .B1(_04474_),
    .B2(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__inv_2 _28416_ (.A(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__o211a_1 _28417_ (.A1(_04464_),
    .A2(net130),
    .B1(net197),
    .C1(_04473_),
    .X(_04478_));
 sky130_fd_sc_hd__o211ai_4 _28418_ (.A1(_04464_),
    .A2(net130),
    .B1(net197),
    .C1(_04473_),
    .Y(_04479_));
 sky130_fd_sc_hd__o221ai_4 _28419_ (.A1(net130),
    .A2(_04465_),
    .B1(_04474_),
    .B2(_04475_),
    .C1(_08313_),
    .Y(_04480_));
 sky130_fd_sc_hd__nand2_1 _28420_ (.A(_04479_),
    .B(_04480_),
    .Y(_04482_));
 sky130_fd_sc_hd__a211oi_1 _28421_ (.A1(_03985_),
    .A2(_03981_),
    .B1(_03803_),
    .C1(_03989_),
    .Y(_04483_));
 sky130_fd_sc_hd__o211a_1 _28422_ (.A1(_04166_),
    .A2(_04174_),
    .B1(_04483_),
    .C1(_04171_),
    .X(_04484_));
 sky130_fd_sc_hd__nand3_1 _28423_ (.A(_04171_),
    .B(_04483_),
    .C(_04176_),
    .Y(_04485_));
 sky130_fd_sc_hd__a31oi_1 _28424_ (.A1(_04344_),
    .A2(_07935_),
    .A3(_04336_),
    .B1(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__a31o_1 _28425_ (.A1(_04344_),
    .A2(_07935_),
    .A3(_04336_),
    .B1(_04485_),
    .X(_04487_));
 sky130_fd_sc_hd__a21oi_1 _28426_ (.A1(_04351_),
    .A2(_04484_),
    .B1(_04352_),
    .Y(_04488_));
 sky130_fd_sc_hd__a211oi_2 _28427_ (.A1(_04347_),
    .A2(_04351_),
    .B1(_04352_),
    .C1(_04486_),
    .Y(_04489_));
 sky130_fd_sc_hd__o211ai_4 _28428_ (.A1(_04348_),
    .A2(_04350_),
    .B1(_04353_),
    .C1(_04487_),
    .Y(_04490_));
 sky130_fd_sc_hd__nand4_4 _28429_ (.A(_04351_),
    .B(_04484_),
    .C(_04353_),
    .D(_03811_),
    .Y(_04491_));
 sky130_fd_sc_hd__nand3_1 _28430_ (.A(_04482_),
    .B(_04490_),
    .C(_04491_),
    .Y(_04493_));
 sky130_fd_sc_hd__a21oi_1 _28431_ (.A1(_04490_),
    .A2(_04491_),
    .B1(_04482_),
    .Y(_04494_));
 sky130_fd_sc_hd__a21o_1 _28432_ (.A1(_04490_),
    .A2(_04491_),
    .B1(_04482_),
    .X(_04495_));
 sky130_fd_sc_hd__o211ai_2 _28433_ (.A1(net137),
    .A2(net134),
    .B1(_04493_),
    .C1(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__or3_1 _28434_ (.A(net137),
    .B(net134),
    .C(_04477_),
    .X(_04497_));
 sky130_fd_sc_hd__a22oi_1 _28435_ (.A1(_04479_),
    .A2(_04480_),
    .B1(_04490_),
    .B2(_04491_),
    .Y(_04498_));
 sky130_fd_sc_hd__a22o_1 _28436_ (.A1(_04479_),
    .A2(_04480_),
    .B1(_04490_),
    .B2(_04491_),
    .X(_04499_));
 sky130_fd_sc_hd__o21ai_2 _28437_ (.A1(net197),
    .A2(_04476_),
    .B1(_04491_),
    .Y(_04500_));
 sky130_fd_sc_hd__a21oi_1 _28438_ (.A1(_04355_),
    .A2(_04488_),
    .B1(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__o211ai_4 _28439_ (.A1(_04476_),
    .A2(net197),
    .B1(_04491_),
    .C1(_04490_),
    .Y(_04502_));
 sky130_fd_sc_hd__a211oi_1 _28440_ (.A1(_04488_),
    .A2(_04355_),
    .B1(_04478_),
    .C1(_04500_),
    .Y(_04505_));
 sky130_fd_sc_hd__o221ai_4 _28441_ (.A1(net137),
    .A2(net134),
    .B1(_04478_),
    .B2(_04502_),
    .C1(_04499_),
    .Y(_04506_));
 sky130_fd_sc_hd__o31a_1 _28442_ (.A1(_10953_),
    .A2(_04498_),
    .A3(_04505_),
    .B1(_04497_),
    .X(_04507_));
 sky130_fd_sc_hd__or3_1 _28443_ (.A(_11459_),
    .B(net129),
    .C(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__o311a_1 _28444_ (.A1(_10953_),
    .A2(_04498_),
    .A3(_04505_),
    .B1(_04497_),
    .C1(_07935_),
    .X(_04509_));
 sky130_fd_sc_hd__o211ai_4 _28445_ (.A1(_10954_),
    .A2(_04477_),
    .B1(_07935_),
    .C1(_04506_),
    .Y(_04510_));
 sky130_fd_sc_hd__o211ai_4 _28446_ (.A1(_04476_),
    .A2(_10954_),
    .B1(_07936_),
    .C1(_04496_),
    .Y(_04511_));
 sky130_fd_sc_hd__a21oi_1 _28447_ (.A1(_07565_),
    .A2(_04362_),
    .B1(_04367_),
    .Y(_04512_));
 sky130_fd_sc_hd__o32a_1 _28448_ (.A1(net221),
    .A2(net219),
    .A3(_04362_),
    .B1(_04363_),
    .B2(_04367_),
    .X(_04513_));
 sky130_fd_sc_hd__a21oi_1 _28449_ (.A1(_04367_),
    .A2(_04365_),
    .B1(_04363_),
    .Y(_04514_));
 sky130_fd_sc_hd__o2bb2ai_1 _28450_ (.A1_N(_04510_),
    .A2_N(_04511_),
    .B1(_04512_),
    .B2(_04366_),
    .Y(_04516_));
 sky130_fd_sc_hd__nand3_1 _28451_ (.A(_04513_),
    .B(_04511_),
    .C(_04510_),
    .Y(_04517_));
 sky130_fd_sc_hd__o211ai_1 _28452_ (.A1(_11459_),
    .A2(net129),
    .B1(_04516_),
    .C1(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__o31a_1 _28453_ (.A1(_11459_),
    .A2(net129),
    .A3(_04507_),
    .B1(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__a21oi_1 _28454_ (.A1(_04508_),
    .A2(_04518_),
    .B1(_07564_),
    .Y(_04520_));
 sky130_fd_sc_hd__a31oi_1 _28455_ (.A1(_11465_),
    .A2(_04516_),
    .A3(_04517_),
    .B1(_07565_),
    .Y(_04521_));
 sky130_fd_sc_hd__o21ai_1 _28456_ (.A1(_11465_),
    .A2(_04507_),
    .B1(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__a21oi_1 _28457_ (.A1(_04508_),
    .A2(_04521_),
    .B1(_04520_),
    .Y(_04523_));
 sky130_fd_sc_hd__o21ai_1 _28458_ (.A1(_04373_),
    .A2(_04375_),
    .B1(_04372_),
    .Y(_04524_));
 sky130_fd_sc_hd__nor2_1 _28459_ (.A(_04523_),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__o21ai_1 _28460_ (.A1(_11944_),
    .A2(_04525_),
    .B1(_04519_),
    .Y(_04527_));
 sky130_fd_sc_hd__nor3b_1 _28461_ (.A(_05051_),
    .B(_04378_),
    .C_N(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__o221a_1 _28462_ (.A1(_04525_),
    .A2(_11944_),
    .B1(_05051_),
    .B2(_04378_),
    .C1(_04519_),
    .X(_04529_));
 sky130_fd_sc_hd__nor2_1 _28463_ (.A(_04528_),
    .B(_04529_),
    .Y(net113));
 sky130_fd_sc_hd__o211a_1 _28464_ (.A1(_11944_),
    .A2(_04525_),
    .B1(_04519_),
    .C1(_04378_),
    .X(_04530_));
 sky130_fd_sc_hd__nor2_1 _28465_ (.A(_05051_),
    .B(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__o211ai_2 _28466_ (.A1(_04380_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_04389_),
    .Y(_04532_));
 sky130_fd_sc_hd__o21ai_4 _28467_ (.A1(net181),
    .A2(net179),
    .B1(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__or3_1 _28468_ (.A(net157),
    .B(_08712_),
    .C(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__and3_1 _28469_ (.A(_04532_),
    .B(net159),
    .C(_10971_),
    .X(_04535_));
 sky130_fd_sc_hd__o2bb2a_1 _28470_ (.A1_N(net159),
    .A2_N(_04532_),
    .B1(_10967_),
    .B2(_10965_),
    .X(_04537_));
 sky130_fd_sc_hd__nor2_1 _28471_ (.A(_04535_),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__o211ai_2 _28472_ (.A1(_04237_),
    .A2(net152),
    .B1(_04395_),
    .C1(_04252_),
    .Y(_04539_));
 sky130_fd_sc_hd__o221ai_4 _28473_ (.A1(_04535_),
    .A2(_04537_),
    .B1(_04397_),
    .B2(_04399_),
    .C1(_04395_),
    .Y(_04540_));
 sky130_fd_sc_hd__o211ai_4 _28474_ (.A1(_10492_),
    .A2(_04391_),
    .B1(_04538_),
    .C1(_04539_),
    .Y(_04541_));
 sky130_fd_sc_hd__nand3_4 _28475_ (.A(_04540_),
    .B(_04541_),
    .C(net149),
    .Y(_04542_));
 sky130_fd_sc_hd__and3_1 _28476_ (.A(_08710_),
    .B(_08713_),
    .C(_04533_),
    .X(_04543_));
 sky130_fd_sc_hd__a21oi_1 _28477_ (.A1(_04540_),
    .A2(_04541_),
    .B1(_08715_),
    .Y(_04544_));
 sky130_fd_sc_hd__o31a_4 _28478_ (.A1(net157),
    .A2(_08712_),
    .A3(_04533_),
    .B1(_04542_),
    .X(_04545_));
 sky130_fd_sc_hd__o21ai_1 _28479_ (.A1(net149),
    .A2(_04533_),
    .B1(_04542_),
    .Y(_04546_));
 sky130_fd_sc_hd__a2bb2oi_1 _28480_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_04534_),
    .B2(_04542_),
    .Y(_04548_));
 sky130_fd_sc_hd__a2bb2o_1 _28481_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_04534_),
    .B2(_04542_),
    .X(_04549_));
 sky130_fd_sc_hd__o211a_2 _28482_ (.A1(net149),
    .A2(_04533_),
    .B1(net150),
    .C1(_04542_),
    .X(_04550_));
 sky130_fd_sc_hd__o211ai_4 _28483_ (.A1(net149),
    .A2(_04533_),
    .B1(net150),
    .C1(_04542_),
    .Y(_04551_));
 sky130_fd_sc_hd__o41ai_2 _28484_ (.A1(net164),
    .A2(_10490_),
    .A3(_04543_),
    .A4(_04544_),
    .B1(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__o2111ai_1 _28485_ (.A1(_04409_),
    .A2(net152),
    .B1(_04549_),
    .C1(_04424_),
    .D1(_04551_),
    .Y(_04553_));
 sky130_fd_sc_hd__o2bb2ai_1 _28486_ (.A1_N(_04412_),
    .A2_N(_04424_),
    .B1(_04548_),
    .B2(_04550_),
    .Y(_04554_));
 sky130_fd_sc_hd__a21oi_4 _28487_ (.A1(_04412_),
    .A2(_04424_),
    .B1(_04552_),
    .Y(_04555_));
 sky130_fd_sc_hd__o211ai_2 _28488_ (.A1(_04548_),
    .A2(_04550_),
    .B1(_04412_),
    .C1(_04424_),
    .Y(_04556_));
 sky130_fd_sc_hd__o211ai_2 _28489_ (.A1(net148),
    .A2(net147),
    .B1(_04553_),
    .C1(_04554_),
    .Y(_04557_));
 sky130_fd_sc_hd__o21ai_4 _28490_ (.A1(net148),
    .A2(net147),
    .B1(_04556_),
    .Y(_04559_));
 sky130_fd_sc_hd__o22ai_4 _28491_ (.A1(net145),
    .A2(_04545_),
    .B1(_04555_),
    .B2(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__inv_2 _28492_ (.A(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__o221ai_4 _28493_ (.A1(net170),
    .A2(net168),
    .B1(_04546_),
    .B2(net145),
    .C1(_04557_),
    .Y(_04562_));
 sky130_fd_sc_hd__inv_2 _28494_ (.A(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__o221a_1 _28495_ (.A1(net145),
    .A2(_04545_),
    .B1(_04555_),
    .B2(_04559_),
    .C1(net152),
    .X(_04564_));
 sky130_fd_sc_hd__o221ai_4 _28496_ (.A1(net145),
    .A2(_04545_),
    .B1(_04555_),
    .B2(_04559_),
    .C1(net152),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _28497_ (.A(_04562_),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__nand4_2 _28498_ (.A(_03933_),
    .B(_03934_),
    .C(_04110_),
    .D(_04112_),
    .Y(_04567_));
 sky130_fd_sc_hd__a211oi_4 _28499_ (.A1(_04262_),
    .A2(_04281_),
    .B1(_04567_),
    .C1(_04286_),
    .Y(_04568_));
 sky130_fd_sc_hd__nand2_1 _28500_ (.A(_04434_),
    .B(_04568_),
    .Y(_04570_));
 sky130_fd_sc_hd__a32oi_1 _28501_ (.A1(net171),
    .A2(_04428_),
    .A3(_04429_),
    .B1(_04434_),
    .B2(_04568_),
    .Y(_04571_));
 sky130_fd_sc_hd__o211ai_4 _28502_ (.A1(_04440_),
    .A2(_04433_),
    .B1(_04435_),
    .C1(_04570_),
    .Y(_04572_));
 sky130_fd_sc_hd__nand3_1 _28503_ (.A(_04434_),
    .B(_04435_),
    .C(_04568_),
    .Y(_04573_));
 sky130_fd_sc_hd__and4_1 _28504_ (.A(_03942_),
    .B(_04434_),
    .C(_04435_),
    .D(_04568_),
    .X(_04574_));
 sky130_fd_sc_hd__nand4_4 _28505_ (.A(_03942_),
    .B(_04434_),
    .C(_04435_),
    .D(_04568_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21oi_2 _28506_ (.A1(_04572_),
    .A2(_04575_),
    .B1(_04566_),
    .Y(_04576_));
 sky130_fd_sc_hd__o211ai_1 _28507_ (.A1(_04573_),
    .A2(_03943_),
    .B1(_04566_),
    .C1(_04572_),
    .Y(_04577_));
 sky130_fd_sc_hd__o21ai_2 _28508_ (.A1(net156),
    .A2(net154),
    .B1(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__a22oi_1 _28509_ (.A1(_04562_),
    .A2(_04565_),
    .B1(_04572_),
    .B2(_04575_),
    .Y(_04579_));
 sky130_fd_sc_hd__a22o_1 _28510_ (.A1(_04562_),
    .A2(_04565_),
    .B1(_04572_),
    .B2(_04575_),
    .X(_04581_));
 sky130_fd_sc_hd__o211ai_4 _28511_ (.A1(_04560_),
    .A2(_10027_),
    .B1(_04575_),
    .C1(_04572_),
    .Y(_04582_));
 sky130_fd_sc_hd__a211oi_1 _28512_ (.A1(_04444_),
    .A2(_04571_),
    .B1(_04566_),
    .C1(_04574_),
    .Y(_04583_));
 sky130_fd_sc_hd__or3_2 _28513_ (.A(net156),
    .B(net154),
    .C(_04561_),
    .X(_04584_));
 sky130_fd_sc_hd__o221ai_4 _28514_ (.A1(net156),
    .A2(net154),
    .B1(_04563_),
    .B2(_04582_),
    .C1(_04581_),
    .Y(_04585_));
 sky130_fd_sc_hd__o22a_1 _28515_ (.A1(net144),
    .A2(_04560_),
    .B1(_04576_),
    .B2(_04578_),
    .X(_04586_));
 sky130_fd_sc_hd__a22o_2 _28516_ (.A1(_09575_),
    .A2(_09577_),
    .B1(_04584_),
    .B2(_04585_),
    .X(_04587_));
 sky130_fd_sc_hd__inv_2 _28517_ (.A(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__o311a_2 _28518_ (.A1(_09562_),
    .A2(_04579_),
    .A3(_04583_),
    .B1(_04584_),
    .C1(_09594_),
    .X(_04589_));
 sky130_fd_sc_hd__nand3_4 _28519_ (.A(_04585_),
    .B(_09594_),
    .C(_04584_),
    .Y(_04590_));
 sky130_fd_sc_hd__o221a_1 _28520_ (.A1(net144),
    .A2(_04560_),
    .B1(_04576_),
    .B2(_04578_),
    .C1(net171),
    .X(_04592_));
 sky130_fd_sc_hd__o221ai_4 _28521_ (.A1(net144),
    .A2(_04560_),
    .B1(_04576_),
    .B2(_04578_),
    .C1(net171),
    .Y(_04593_));
 sky130_fd_sc_hd__o211a_1 _28522_ (.A1(net176),
    .A2(_04297_),
    .B1(_04450_),
    .C1(_04454_),
    .X(_04594_));
 sky130_fd_sc_hd__o211ai_2 _28523_ (.A1(net176),
    .A2(_04297_),
    .B1(_04450_),
    .C1(_04454_),
    .Y(_04595_));
 sky130_fd_sc_hd__o21ai_4 _28524_ (.A1(_09139_),
    .A2(_04447_),
    .B1(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__a21oi_4 _28525_ (.A1(_04590_),
    .A2(_04593_),
    .B1(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__a21o_1 _28526_ (.A1(_04590_),
    .A2(_04593_),
    .B1(_04596_),
    .X(_04598_));
 sky130_fd_sc_hd__o211a_1 _28527_ (.A1(_04455_),
    .A2(_04594_),
    .B1(_04593_),
    .C1(_04590_),
    .X(_04599_));
 sky130_fd_sc_hd__nand3_2 _28528_ (.A(_04590_),
    .B(_04596_),
    .C(_04593_),
    .Y(_04600_));
 sky130_fd_sc_hd__a31oi_2 _28529_ (.A1(_04590_),
    .A2(_04596_),
    .A3(_04593_),
    .B1(_09578_),
    .Y(_04601_));
 sky130_fd_sc_hd__a31o_1 _28530_ (.A1(_04590_),
    .A2(_04596_),
    .A3(_04593_),
    .B1(_09578_),
    .X(_04603_));
 sky130_fd_sc_hd__nand2_1 _28531_ (.A(_04601_),
    .B(_04598_),
    .Y(_04604_));
 sky130_fd_sc_hd__o22ai_2 _28532_ (.A1(net142),
    .A2(_09573_),
    .B1(_04597_),
    .B2(_04599_),
    .Y(_04605_));
 sky130_fd_sc_hd__a21oi_4 _28533_ (.A1(_04601_),
    .A2(_04598_),
    .B1(_04588_),
    .Y(_04606_));
 sky130_fd_sc_hd__a31o_2 _28534_ (.A1(net132),
    .A2(_04598_),
    .A3(_04600_),
    .B1(_04588_),
    .X(_04607_));
 sky130_fd_sc_hd__o211ai_4 _28535_ (.A1(_04340_),
    .A2(_04328_),
    .B1(_04315_),
    .C1(_04466_),
    .Y(_04608_));
 sky130_fd_sc_hd__a31oi_2 _28536_ (.A1(_04315_),
    .A2(_04342_),
    .A3(_04466_),
    .B1(_04467_),
    .Y(_04609_));
 sky130_fd_sc_hd__o21ai_2 _28537_ (.A1(_04597_),
    .A2(_04603_),
    .B1(_09139_),
    .Y(_04610_));
 sky130_fd_sc_hd__o211a_1 _28538_ (.A1(_04597_),
    .A2(_04603_),
    .B1(_09139_),
    .C1(_04587_),
    .X(_04611_));
 sky130_fd_sc_hd__o211ai_4 _28539_ (.A1(_04597_),
    .A2(_04603_),
    .B1(_09139_),
    .C1(_04587_),
    .Y(_04612_));
 sky130_fd_sc_hd__a2bb2oi_4 _28540_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_04587_),
    .B2(_04604_),
    .Y(_04615_));
 sky130_fd_sc_hd__o221ai_4 _28541_ (.A1(net194),
    .A2(net190),
    .B1(net132),
    .B2(_04586_),
    .C1(_04605_),
    .Y(_04616_));
 sky130_fd_sc_hd__o21ai_1 _28542_ (.A1(_04588_),
    .A2(_04610_),
    .B1(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__o2111a_1 _28543_ (.A1(_04469_),
    .A2(_04471_),
    .B1(_04612_),
    .C1(_04616_),
    .D1(_04466_),
    .X(_04618_));
 sky130_fd_sc_hd__a2bb2o_2 _28544_ (.A1_N(net141),
    .A2_N(net139),
    .B1(_04609_),
    .B2(_04617_),
    .X(_04619_));
 sky130_fd_sc_hd__o221ai_4 _28545_ (.A1(_04464_),
    .A2(net176),
    .B1(_09139_),
    .B2(_04606_),
    .C1(_04608_),
    .Y(_04620_));
 sky130_fd_sc_hd__o2bb2ai_1 _28546_ (.A1_N(_04468_),
    .A2_N(_04608_),
    .B1(_04611_),
    .B2(_04615_),
    .Y(_04621_));
 sky130_fd_sc_hd__or3_1 _28547_ (.A(net141),
    .B(net139),
    .C(_04606_),
    .X(_04622_));
 sky130_fd_sc_hd__o221ai_4 _28548_ (.A1(net141),
    .A2(net139),
    .B1(_04611_),
    .B2(_04620_),
    .C1(_04621_),
    .Y(_04623_));
 sky130_fd_sc_hd__o22a_4 _28549_ (.A1(net130),
    .A2(_04607_),
    .B1(_04618_),
    .B2(_04619_),
    .X(_04624_));
 sky130_fd_sc_hd__and3_1 _28550_ (.A(_04623_),
    .B(net178),
    .C(_04622_),
    .X(_04626_));
 sky130_fd_sc_hd__o211ai_2 _28551_ (.A1(net130),
    .A2(_04606_),
    .B1(net178),
    .C1(_04623_),
    .Y(_04627_));
 sky130_fd_sc_hd__a2bb2oi_2 _28552_ (.A1_N(_08724_),
    .A2_N(net196),
    .B1(_04622_),
    .B2(_04623_),
    .Y(_04628_));
 sky130_fd_sc_hd__o221ai_4 _28553_ (.A1(net130),
    .A2(_04607_),
    .B1(_04618_),
    .B2(_04619_),
    .C1(net176),
    .Y(_04629_));
 sky130_fd_sc_hd__nor2_1 _28554_ (.A(_04626_),
    .B(_04628_),
    .Y(_04630_));
 sky130_fd_sc_hd__o2bb2ai_1 _28555_ (.A1_N(_04479_),
    .A2_N(_04502_),
    .B1(_04626_),
    .B2(_04628_),
    .Y(_04631_));
 sky130_fd_sc_hd__o2111ai_4 _28556_ (.A1(_04477_),
    .A2(_08313_),
    .B1(_04627_),
    .C1(_04502_),
    .D1(_04629_),
    .Y(_04632_));
 sky130_fd_sc_hd__o211ai_1 _28557_ (.A1(_04478_),
    .A2(_04501_),
    .B1(_04627_),
    .C1(_04629_),
    .Y(_04633_));
 sky130_fd_sc_hd__o221ai_2 _28558_ (.A1(_04477_),
    .A2(_08313_),
    .B1(_04628_),
    .B2(_04626_),
    .C1(_04502_),
    .Y(_04634_));
 sky130_fd_sc_hd__a22oi_4 _28559_ (.A1(_10950_),
    .A2(_10952_),
    .B1(_04631_),
    .B2(_04632_),
    .Y(_04635_));
 sky130_fd_sc_hd__o211ai_1 _28560_ (.A1(net137),
    .A2(net134),
    .B1(_04633_),
    .C1(_04634_),
    .Y(_04637_));
 sky130_fd_sc_hd__o221a_1 _28561_ (.A1(net130),
    .A2(_04607_),
    .B1(_04618_),
    .B2(_04619_),
    .C1(_10953_),
    .X(_04638_));
 sky130_fd_sc_hd__a21oi_4 _28562_ (.A1(_10953_),
    .A2(_04624_),
    .B1(_04635_),
    .Y(_04639_));
 sky130_fd_sc_hd__o22a_1 _28563_ (.A1(_08307_),
    .A2(net216),
    .B1(_04635_),
    .B2(_04638_),
    .X(_04640_));
 sky130_fd_sc_hd__o21ai_1 _28564_ (.A1(_04635_),
    .A2(_04638_),
    .B1(net197),
    .Y(_04641_));
 sky130_fd_sc_hd__a31o_1 _28565_ (.A1(_10954_),
    .A2(_04633_),
    .A3(_04634_),
    .B1(net197),
    .X(_04642_));
 sky130_fd_sc_hd__nand3b_2 _28566_ (.A_N(_04638_),
    .B(_08313_),
    .C(_04637_),
    .Y(_04643_));
 sky130_fd_sc_hd__o2111a_1 _28567_ (.A1(_04000_),
    .A2(_03995_),
    .B1(_03999_),
    .C1(_04189_),
    .D1(_04191_),
    .X(_04644_));
 sky130_fd_sc_hd__and3_1 _28568_ (.A(_04364_),
    .B(_04644_),
    .C(_04365_),
    .X(_04645_));
 sky130_fd_sc_hd__nand3_1 _28569_ (.A(_04364_),
    .B(_04644_),
    .C(_04365_),
    .Y(_04646_));
 sky130_fd_sc_hd__a31o_1 _28570_ (.A1(_04506_),
    .A2(_07935_),
    .A3(_04497_),
    .B1(_04646_),
    .X(_04648_));
 sky130_fd_sc_hd__o211a_1 _28571_ (.A1(_04514_),
    .A2(_04509_),
    .B1(_04511_),
    .C1(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__o211ai_2 _28572_ (.A1(_04514_),
    .A2(_04509_),
    .B1(_04511_),
    .C1(_04648_),
    .Y(_04650_));
 sky130_fd_sc_hd__nand4_4 _28573_ (.A(_04645_),
    .B(_04511_),
    .C(_04510_),
    .D(_04011_),
    .Y(_04651_));
 sky130_fd_sc_hd__a41o_1 _28574_ (.A1(_04011_),
    .A2(_04510_),
    .A3(_04511_),
    .A4(_04645_),
    .B1(_04649_),
    .X(_04652_));
 sky130_fd_sc_hd__a22o_1 _28575_ (.A1(_04641_),
    .A2(_04643_),
    .B1(_04650_),
    .B2(_04651_),
    .X(_04653_));
 sky130_fd_sc_hd__o31ai_1 _28576_ (.A1(net197),
    .A2(_04635_),
    .A3(_04638_),
    .B1(_04651_),
    .Y(_04654_));
 sky130_fd_sc_hd__nand3_4 _28577_ (.A(_04643_),
    .B(_04650_),
    .C(_04651_),
    .Y(_04655_));
 sky130_fd_sc_hd__o221ai_4 _28578_ (.A1(_11459_),
    .A2(net129),
    .B1(_04640_),
    .B2(_04655_),
    .C1(_04653_),
    .Y(_04656_));
 sky130_fd_sc_hd__o21ai_1 _28579_ (.A1(_11465_),
    .A2(_04639_),
    .B1(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__o311a_1 _28580_ (.A1(_11459_),
    .A2(net129),
    .A3(_04639_),
    .B1(_07935_),
    .C1(_04656_),
    .X(_04659_));
 sky130_fd_sc_hd__o211ai_2 _28581_ (.A1(_11465_),
    .A2(_04639_),
    .B1(_07935_),
    .C1(_04656_),
    .Y(_04660_));
 sky130_fd_sc_hd__o21ai_2 _28582_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_04657_),
    .Y(_04661_));
 sky130_fd_sc_hd__a21oi_1 _28583_ (.A1(_04524_),
    .A2(_04522_),
    .B1(_04520_),
    .Y(_04662_));
 sky130_fd_sc_hd__a221oi_1 _28584_ (.A1(_04524_),
    .A2(_04522_),
    .B1(_04661_),
    .B2(_04660_),
    .C1(_04520_),
    .Y(_04663_));
 sky130_fd_sc_hd__o221a_1 _28585_ (.A1(_11465_),
    .A2(_04639_),
    .B1(_11944_),
    .B2(_04663_),
    .C1(_04656_),
    .X(_04664_));
 sky130_fd_sc_hd__xnor2_1 _28586_ (.A(_04531_),
    .B(_04664_),
    .Y(net114));
 sky130_fd_sc_hd__nand2_1 _28587_ (.A(_04530_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__a2bb2o_1 _28588_ (.A1_N(_04832_),
    .A2_N(_04942_),
    .B1(_04530_),
    .B2(_04664_),
    .X(_04666_));
 sky130_fd_sc_hd__o211ai_4 _28589_ (.A1(_04533_),
    .A2(_10970_),
    .B1(_11471_),
    .C1(_04541_),
    .Y(_04667_));
 sky130_fd_sc_hd__o21ai_2 _28590_ (.A1(net157),
    .A2(_08712_),
    .B1(_04667_),
    .Y(_04669_));
 sky130_fd_sc_hd__inv_2 _28591_ (.A(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__and3_1 _28592_ (.A(_04667_),
    .B(net149),
    .C(_10971_),
    .X(_04671_));
 sky130_fd_sc_hd__o211ai_4 _28593_ (.A1(net157),
    .A2(_08712_),
    .B1(_10971_),
    .C1(_04667_),
    .Y(_04672_));
 sky130_fd_sc_hd__a31o_1 _28594_ (.A1(_08706_),
    .A2(_08708_),
    .A3(_04667_),
    .B1(_10971_),
    .X(_04673_));
 sky130_fd_sc_hd__and2_1 _28595_ (.A(_04672_),
    .B(_04673_),
    .X(_04674_));
 sky130_fd_sc_hd__nand2_1 _28596_ (.A(_04672_),
    .B(_04673_),
    .Y(_04675_));
 sky130_fd_sc_hd__o221ai_4 _28597_ (.A1(net152),
    .A2(_04409_),
    .B1(_04545_),
    .B2(_10491_),
    .C1(_04424_),
    .Y(_04676_));
 sky130_fd_sc_hd__a31oi_1 _28598_ (.A1(_04412_),
    .A2(_04424_),
    .A3(_04549_),
    .B1(_04550_),
    .Y(_04677_));
 sky130_fd_sc_hd__a311oi_4 _28599_ (.A1(_04412_),
    .A2(_04424_),
    .A3(_04549_),
    .B1(_04550_),
    .C1(_04675_),
    .Y(_04678_));
 sky130_fd_sc_hd__nand4_2 _28600_ (.A(_04551_),
    .B(_04672_),
    .C(_04673_),
    .D(_04676_),
    .Y(_04680_));
 sky130_fd_sc_hd__a21oi_1 _28601_ (.A1(_04551_),
    .A2(_04676_),
    .B1(_04674_),
    .Y(_04681_));
 sky130_fd_sc_hd__o211ai_2 _28602_ (.A1(_04674_),
    .A2(_04677_),
    .B1(_04680_),
    .C1(net145),
    .Y(_04682_));
 sky130_fd_sc_hd__o22ai_4 _28603_ (.A1(net148),
    .A2(net147),
    .B1(_04678_),
    .B2(_04681_),
    .Y(_04683_));
 sky130_fd_sc_hd__o21a_2 _28604_ (.A1(net145),
    .A2(_04669_),
    .B1(_04682_),
    .X(_04684_));
 sky130_fd_sc_hd__o221a_2 _28605_ (.A1(_09559_),
    .A2(_09560_),
    .B1(_04670_),
    .B2(net145),
    .C1(_04683_),
    .X(_04685_));
 sky130_fd_sc_hd__o211a_1 _28606_ (.A1(_04670_),
    .A2(net145),
    .B1(_10492_),
    .C1(_04683_),
    .X(_04686_));
 sky130_fd_sc_hd__o211ai_4 _28607_ (.A1(_04670_),
    .A2(net145),
    .B1(_10492_),
    .C1(_04683_),
    .Y(_04687_));
 sky130_fd_sc_hd__o211ai_4 _28608_ (.A1(net145),
    .A2(_04669_),
    .B1(_10491_),
    .C1(_04682_),
    .Y(_04688_));
 sky130_fd_sc_hd__nand2_2 _28609_ (.A(_04687_),
    .B(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__a21oi_1 _28610_ (.A1(_04572_),
    .A2(_04575_),
    .B1(_04563_),
    .Y(_04691_));
 sky130_fd_sc_hd__o2bb2ai_1 _28611_ (.A1_N(_04572_),
    .A2_N(_04575_),
    .B1(net152),
    .B2(_04561_),
    .Y(_04692_));
 sky130_fd_sc_hd__a21oi_4 _28612_ (.A1(_04562_),
    .A2(_04582_),
    .B1(_04689_),
    .Y(_04693_));
 sky130_fd_sc_hd__o2111ai_4 _28613_ (.A1(_10027_),
    .A2(_04560_),
    .B1(_04687_),
    .C1(_04688_),
    .D1(_04692_),
    .Y(_04694_));
 sky130_fd_sc_hd__o211ai_1 _28614_ (.A1(net152),
    .A2(_04561_),
    .B1(_04582_),
    .C1(_04689_),
    .Y(_04695_));
 sky130_fd_sc_hd__a31o_1 _28615_ (.A1(_04562_),
    .A2(_04582_),
    .A3(_04689_),
    .B1(_09562_),
    .X(_04696_));
 sky130_fd_sc_hd__o311a_2 _28616_ (.A1(_04564_),
    .A2(_04689_),
    .A3(_04691_),
    .B1(_04695_),
    .C1(net144),
    .X(_04697_));
 sky130_fd_sc_hd__o22a_1 _28617_ (.A1(net144),
    .A2(_04684_),
    .B1(_04693_),
    .B2(_04696_),
    .X(_04698_));
 sky130_fd_sc_hd__o211a_1 _28618_ (.A1(_04685_),
    .A2(_04697_),
    .B1(_09572_),
    .C1(_09574_),
    .X(_04699_));
 sky130_fd_sc_hd__or3_4 _28619_ (.A(net142),
    .B(_09573_),
    .C(_04698_),
    .X(_04700_));
 sky130_fd_sc_hd__o22a_1 _28620_ (.A1(net170),
    .A2(net168),
    .B1(_04685_),
    .B2(_04697_),
    .X(_04702_));
 sky130_fd_sc_hd__o22ai_4 _28621_ (.A1(net170),
    .A2(net168),
    .B1(_04685_),
    .B2(_04697_),
    .Y(_04703_));
 sky130_fd_sc_hd__o221ai_4 _28622_ (.A1(net144),
    .A2(_04684_),
    .B1(_04693_),
    .B2(_04696_),
    .C1(net152),
    .Y(_04704_));
 sky130_fd_sc_hd__nand2_1 _28623_ (.A(_04703_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__nand4_1 _28624_ (.A(_04130_),
    .B(_04131_),
    .C(_04299_),
    .D(_04300_),
    .Y(_04706_));
 sky130_fd_sc_hd__a211oi_2 _28625_ (.A1(_04432_),
    .A2(_04452_),
    .B1(_04706_),
    .C1(_04455_),
    .Y(_04707_));
 sky130_fd_sc_hd__nand4_4 _28626_ (.A(_04456_),
    .B(_04301_),
    .C(_04132_),
    .D(_04454_),
    .Y(_04708_));
 sky130_fd_sc_hd__a31oi_2 _28627_ (.A1(_04585_),
    .A2(_09594_),
    .A3(_04584_),
    .B1(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__a211oi_4 _28628_ (.A1(_04596_),
    .A2(_04590_),
    .B1(_04592_),
    .C1(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__o211ai_4 _28629_ (.A1(_04708_),
    .A2(_04589_),
    .B1(_04593_),
    .C1(_04600_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand3_2 _28630_ (.A(_04707_),
    .B(_04593_),
    .C(_04141_),
    .Y(_04713_));
 sky130_fd_sc_hd__nand4_4 _28631_ (.A(_04590_),
    .B(_04707_),
    .C(_04593_),
    .D(_04141_),
    .Y(_04714_));
 sky130_fd_sc_hd__o211ai_2 _28632_ (.A1(_04589_),
    .A2(_04713_),
    .B1(_04711_),
    .C1(_04705_),
    .Y(_04715_));
 sky130_fd_sc_hd__a21o_1 _28633_ (.A1(_04711_),
    .A2(_04714_),
    .B1(_04705_),
    .X(_04716_));
 sky130_fd_sc_hd__a22o_2 _28634_ (.A1(_04703_),
    .A2(_04704_),
    .B1(_04711_),
    .B2(_04714_),
    .X(_04717_));
 sky130_fd_sc_hd__nand2_1 _28635_ (.A(_04704_),
    .B(_04714_),
    .Y(_04718_));
 sky130_fd_sc_hd__o211ai_4 _28636_ (.A1(_04713_),
    .A2(_04589_),
    .B1(_04704_),
    .C1(_04711_),
    .Y(_04719_));
 sky130_fd_sc_hd__nand4_2 _28637_ (.A(_04703_),
    .B(_04704_),
    .C(_04711_),
    .D(_04714_),
    .Y(_04720_));
 sky130_fd_sc_hd__o221ai_4 _28638_ (.A1(net142),
    .A2(_09573_),
    .B1(_04702_),
    .B2(_04719_),
    .C1(_04717_),
    .Y(_04721_));
 sky130_fd_sc_hd__or4_2 _28639_ (.A(net142),
    .B(_09573_),
    .C(_04685_),
    .D(_04697_),
    .X(_04722_));
 sky130_fd_sc_hd__o211ai_4 _28640_ (.A1(net142),
    .A2(_09573_),
    .B1(_04715_),
    .C1(_04716_),
    .Y(_04724_));
 sky130_fd_sc_hd__a31o_1 _28641_ (.A1(net132),
    .A2(_04717_),
    .A3(_04720_),
    .B1(_04699_),
    .X(_04725_));
 sky130_fd_sc_hd__o311a_2 _28642_ (.A1(net132),
    .A2(_04685_),
    .A3(_04697_),
    .B1(_10479_),
    .C1(_04724_),
    .X(_04726_));
 sky130_fd_sc_hd__a211o_1 _28643_ (.A1(_04700_),
    .A2(_04721_),
    .B1(net141),
    .C1(net139),
    .X(_04727_));
 sky130_fd_sc_hd__a311oi_4 _28644_ (.A1(net132),
    .A2(_04717_),
    .A3(_04720_),
    .B1(net171),
    .C1(_04699_),
    .Y(_04728_));
 sky130_fd_sc_hd__nand3_4 _28645_ (.A(_04721_),
    .B(_09594_),
    .C(_04700_),
    .Y(_04729_));
 sky130_fd_sc_hd__a2bb2oi_1 _28646_ (.A1_N(net189),
    .A2_N(net186),
    .B1(_04700_),
    .B2(_04721_),
    .Y(_04730_));
 sky130_fd_sc_hd__o211ai_4 _28647_ (.A1(net189),
    .A2(net186),
    .B1(_04722_),
    .C1(_04724_),
    .Y(_04731_));
 sky130_fd_sc_hd__o221a_1 _28648_ (.A1(_09139_),
    .A2(_04606_),
    .B1(_04467_),
    .B2(_04471_),
    .C1(_04466_),
    .X(_04732_));
 sky130_fd_sc_hd__o211a_1 _28649_ (.A1(_04464_),
    .A2(net176),
    .B1(_04612_),
    .C1(_04608_),
    .X(_04733_));
 sky130_fd_sc_hd__a31o_1 _28650_ (.A1(_04468_),
    .A2(_04608_),
    .A3(_04612_),
    .B1(_04615_),
    .X(_04735_));
 sky130_fd_sc_hd__a21oi_2 _28651_ (.A1(_04609_),
    .A2(_04612_),
    .B1(_04615_),
    .Y(_04736_));
 sky130_fd_sc_hd__a21oi_1 _28652_ (.A1(_04729_),
    .A2(_04731_),
    .B1(_04735_),
    .Y(_04737_));
 sky130_fd_sc_hd__o2bb2ai_2 _28653_ (.A1_N(_04729_),
    .A2_N(_04731_),
    .B1(_04732_),
    .B2(_04611_),
    .Y(_04738_));
 sky130_fd_sc_hd__o211a_1 _28654_ (.A1(_04615_),
    .A2(_04733_),
    .B1(_04731_),
    .C1(_04729_),
    .X(_04739_));
 sky130_fd_sc_hd__o211ai_4 _28655_ (.A1(_04615_),
    .A2(_04733_),
    .B1(_04731_),
    .C1(_04729_),
    .Y(_04740_));
 sky130_fd_sc_hd__o211ai_2 _28656_ (.A1(net141),
    .A2(net139),
    .B1(_04738_),
    .C1(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__o22ai_2 _28657_ (.A1(net141),
    .A2(net139),
    .B1(_04737_),
    .B2(_04739_),
    .Y(_04742_));
 sky130_fd_sc_hd__o31a_2 _28658_ (.A1(_10479_),
    .A2(_04737_),
    .A3(_04739_),
    .B1(_04727_),
    .X(_04743_));
 sky130_fd_sc_hd__a311o_2 _28659_ (.A1(net130),
    .A2(_04738_),
    .A3(_04740_),
    .B1(_10954_),
    .C1(_04726_),
    .X(_04744_));
 sky130_fd_sc_hd__a2bb2oi_2 _28660_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_04727_),
    .B2(_04741_),
    .Y(_04746_));
 sky130_fd_sc_hd__o221ai_4 _28661_ (.A1(net194),
    .A2(net190),
    .B1(net130),
    .B2(_04725_),
    .C1(_04742_),
    .Y(_04747_));
 sky130_fd_sc_hd__a31o_1 _28662_ (.A1(net130),
    .A2(_04738_),
    .A3(_04740_),
    .B1(_09140_),
    .X(_04748_));
 sky130_fd_sc_hd__a311oi_4 _28663_ (.A1(net130),
    .A2(_04738_),
    .A3(_04740_),
    .B1(_04726_),
    .C1(_09140_),
    .Y(_04749_));
 sky130_fd_sc_hd__nand3_2 _28664_ (.A(_04741_),
    .B(_09139_),
    .C(_04727_),
    .Y(_04750_));
 sky130_fd_sc_hd__o211ai_4 _28665_ (.A1(_04500_),
    .A2(_04489_),
    .B1(_04479_),
    .C1(_04629_),
    .Y(_04751_));
 sky130_fd_sc_hd__o21ai_1 _28666_ (.A1(net176),
    .A2(_04624_),
    .B1(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__o211ai_2 _28667_ (.A1(_04748_),
    .A2(_04726_),
    .B1(_04747_),
    .C1(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__o221ai_4 _28668_ (.A1(_04624_),
    .A2(net176),
    .B1(_04749_),
    .B2(_04746_),
    .C1(_04751_),
    .Y(_04754_));
 sky130_fd_sc_hd__o211ai_4 _28669_ (.A1(net137),
    .A2(net134),
    .B1(_04753_),
    .C1(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__o21ai_1 _28670_ (.A1(_04746_),
    .A2(_04749_),
    .B1(_04752_),
    .Y(_04757_));
 sky130_fd_sc_hd__o2111ai_1 _28671_ (.A1(_04624_),
    .A2(net176),
    .B1(_04750_),
    .C1(_04747_),
    .D1(_04751_),
    .Y(_04758_));
 sky130_fd_sc_hd__o211ai_2 _28672_ (.A1(net137),
    .A2(net134),
    .B1(_04757_),
    .C1(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__o21ai_1 _28673_ (.A1(_10954_),
    .A2(_04743_),
    .B1(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__nand2_2 _28674_ (.A(_04744_),
    .B(_04755_),
    .Y(_04761_));
 sky130_fd_sc_hd__o22ai_1 _28675_ (.A1(_08313_),
    .A2(_04639_),
    .B1(_04654_),
    .B2(_04649_),
    .Y(_04762_));
 sky130_fd_sc_hd__o211ai_4 _28676_ (.A1(_10954_),
    .A2(_04743_),
    .B1(_08730_),
    .C1(_04759_),
    .Y(_04763_));
 sky130_fd_sc_hd__o211ai_4 _28677_ (.A1(_08724_),
    .A2(net196),
    .B1(_04744_),
    .C1(_04755_),
    .Y(_04764_));
 sky130_fd_sc_hd__nand2_1 _28678_ (.A(_04763_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__o2111ai_4 _28679_ (.A1(_08313_),
    .A2(_04639_),
    .B1(_04655_),
    .C1(_04763_),
    .D1(_04764_),
    .Y(_04766_));
 sky130_fd_sc_hd__a21oi_2 _28680_ (.A1(_04762_),
    .A2(_04765_),
    .B1(_11464_),
    .Y(_04768_));
 sky130_fd_sc_hd__a22oi_4 _28681_ (.A1(_11464_),
    .A2(_04761_),
    .B1(_04768_),
    .B2(_04766_),
    .Y(_04769_));
 sky130_fd_sc_hd__a221o_1 _28682_ (.A1(_11464_),
    .A2(_04761_),
    .B1(_04768_),
    .B2(_04766_),
    .C1(_08313_),
    .X(_04770_));
 sky130_fd_sc_hd__xor2_1 _28683_ (.A(net197),
    .B(_04769_),
    .X(_04771_));
 sky130_fd_sc_hd__xor2_1 _28684_ (.A(_08313_),
    .B(_04769_),
    .X(_04772_));
 sky130_fd_sc_hd__and3_1 _28685_ (.A(_04372_),
    .B(_04374_),
    .C(_04205_),
    .X(_04773_));
 sky130_fd_sc_hd__nand3_1 _28686_ (.A(_04660_),
    .B(_04773_),
    .C(_04523_),
    .Y(_04774_));
 sky130_fd_sc_hd__o211ai_2 _28687_ (.A1(_04662_),
    .A2(_04659_),
    .B1(_04661_),
    .C1(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__nand4b_1 _28688_ (.A_N(_04520_),
    .B(_04773_),
    .C(_04522_),
    .D(_04202_),
    .Y(_04776_));
 sky130_fd_sc_hd__nand3b_1 _28689_ (.A_N(_04776_),
    .B(_04661_),
    .C(_04660_),
    .Y(_04777_));
 sky130_fd_sc_hd__nand2_1 _28690_ (.A(_04775_),
    .B(_04777_),
    .Y(_04779_));
 sky130_fd_sc_hd__o211ai_2 _28691_ (.A1(_04769_),
    .A2(net197),
    .B1(_04777_),
    .C1(_04775_),
    .Y(_04780_));
 sky130_fd_sc_hd__a21o_1 _28692_ (.A1(net197),
    .A2(_04769_),
    .B1(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__nand2_1 _28693_ (.A(_04772_),
    .B(_04779_),
    .Y(_04782_));
 sky130_fd_sc_hd__a31o_1 _28694_ (.A1(_04781_),
    .A2(_04782_),
    .A3(net133),
    .B1(_04769_),
    .X(_04783_));
 sky130_fd_sc_hd__xnor2_1 _28695_ (.A(_04666_),
    .B(_04783_),
    .Y(net115));
 sky130_fd_sc_hd__nor2_1 _28696_ (.A(_04665_),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__a31o_1 _28697_ (.A1(_11471_),
    .A2(_04672_),
    .A3(_04680_),
    .B1(_09124_),
    .X(_04785_));
 sky130_fd_sc_hd__o311a_2 _28698_ (.A1(_11470_),
    .A2(_04671_),
    .A3(_04678_),
    .B1(_09562_),
    .C1(net145),
    .X(_04786_));
 sky130_fd_sc_hd__a311o_1 _28699_ (.A1(_11471_),
    .A2(_04672_),
    .A3(_04680_),
    .B1(net144),
    .C1(_09124_),
    .X(_04787_));
 sky130_fd_sc_hd__o311a_1 _28700_ (.A1(_11470_),
    .A2(_04671_),
    .A3(_04678_),
    .B1(_10971_),
    .C1(net145),
    .X(_04789_));
 sky130_fd_sc_hd__and3_1 _28701_ (.A(_10963_),
    .B(_10964_),
    .C(_04785_),
    .X(_04790_));
 sky130_fd_sc_hd__nor2_1 _28702_ (.A(_04789_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__o21a_1 _28703_ (.A1(_04686_),
    .A2(_04693_),
    .B1(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__o21ai_4 _28704_ (.A1(_04686_),
    .A2(_04693_),
    .B1(_04791_),
    .Y(_04793_));
 sky130_fd_sc_hd__o221ai_4 _28705_ (.A1(_10491_),
    .A2(_04684_),
    .B1(_04789_),
    .B2(_04790_),
    .C1(_04694_),
    .Y(_04794_));
 sky130_fd_sc_hd__o211ai_2 _28706_ (.A1(net156),
    .A2(net154),
    .B1(_04793_),
    .C1(_04794_),
    .Y(_04795_));
 sky130_fd_sc_hd__a31o_1 _28707_ (.A1(net144),
    .A2(_04793_),
    .A3(_04794_),
    .B1(_04786_),
    .X(_04796_));
 sky130_fd_sc_hd__o311a_1 _28708_ (.A1(net156),
    .A2(net154),
    .A3(_04785_),
    .B1(_09578_),
    .C1(_04795_),
    .X(_04797_));
 sky130_fd_sc_hd__a311o_1 _28709_ (.A1(net144),
    .A2(_04793_),
    .A3(_04794_),
    .B1(net132),
    .C1(_04786_),
    .X(_04798_));
 sky130_fd_sc_hd__a2bb2oi_1 _28710_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_04787_),
    .B2(_04795_),
    .Y(_04800_));
 sky130_fd_sc_hd__o21ai_2 _28711_ (.A1(_10487_),
    .A2(net165),
    .B1(_04796_),
    .Y(_04801_));
 sky130_fd_sc_hd__a311oi_4 _28712_ (.A1(net144),
    .A2(_04793_),
    .A3(_04794_),
    .B1(_10492_),
    .C1(_04786_),
    .Y(_04802_));
 sky130_fd_sc_hd__a311o_1 _28713_ (.A1(net144),
    .A2(_04793_),
    .A3(_04794_),
    .B1(_10492_),
    .C1(_04786_),
    .X(_04803_));
 sky130_fd_sc_hd__o22ai_1 _28714_ (.A1(net152),
    .A2(_04698_),
    .B1(_04718_),
    .B2(_04710_),
    .Y(_04804_));
 sky130_fd_sc_hd__a31oi_1 _28715_ (.A1(_04704_),
    .A2(_04711_),
    .A3(_04714_),
    .B1(_04702_),
    .Y(_04805_));
 sky130_fd_sc_hd__o2111ai_4 _28716_ (.A1(_04718_),
    .A2(_04710_),
    .B1(_04703_),
    .C1(_04803_),
    .D1(_04801_),
    .Y(_04806_));
 sky130_fd_sc_hd__o2bb2ai_2 _28717_ (.A1_N(_04703_),
    .A2_N(_04719_),
    .B1(_04800_),
    .B2(_04802_),
    .Y(_04807_));
 sky130_fd_sc_hd__o211ai_2 _28718_ (.A1(net142),
    .A2(_09573_),
    .B1(_04806_),
    .C1(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__a22o_1 _28719_ (.A1(_09575_),
    .A2(_09577_),
    .B1(_04787_),
    .B2(_04795_),
    .X(_04809_));
 sky130_fd_sc_hd__nand3_1 _28720_ (.A(_04804_),
    .B(_04803_),
    .C(_04801_),
    .Y(_04811_));
 sky130_fd_sc_hd__o221ai_1 _28721_ (.A1(_04718_),
    .A2(_04710_),
    .B1(_04802_),
    .B2(_04800_),
    .C1(_04703_),
    .Y(_04812_));
 sky130_fd_sc_hd__o211ai_1 _28722_ (.A1(net142),
    .A2(_09573_),
    .B1(_04811_),
    .C1(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__a31oi_4 _28723_ (.A1(net132),
    .A2(_04806_),
    .A3(_04807_),
    .B1(_04797_),
    .Y(_04814_));
 sky130_fd_sc_hd__a31o_1 _28724_ (.A1(net132),
    .A2(_04806_),
    .A3(_04807_),
    .B1(_04797_),
    .X(_04815_));
 sky130_fd_sc_hd__and3_1 _28725_ (.A(_10027_),
    .B(_04798_),
    .C(_04808_),
    .X(_04816_));
 sky130_fd_sc_hd__o211ai_4 _28726_ (.A1(net170),
    .A2(net168),
    .B1(_04798_),
    .C1(_04808_),
    .Y(_04817_));
 sky130_fd_sc_hd__and3_1 _28727_ (.A(_04813_),
    .B(net152),
    .C(_04809_),
    .X(_04818_));
 sky130_fd_sc_hd__nand3_1 _28728_ (.A(_04813_),
    .B(net152),
    .C(_04809_),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_1 _28729_ (.A(_04817_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__and3_1 _28730_ (.A(_04320_),
    .B(_04466_),
    .C(_04468_),
    .X(_04822_));
 sky130_fd_sc_hd__o211a_1 _28731_ (.A1(_04588_),
    .A2(_04610_),
    .B1(_04822_),
    .C1(_04616_),
    .X(_04823_));
 sky130_fd_sc_hd__o211ai_2 _28732_ (.A1(_04588_),
    .A2(_04610_),
    .B1(_04822_),
    .C1(_04616_),
    .Y(_04824_));
 sky130_fd_sc_hd__a31oi_2 _28733_ (.A1(_04721_),
    .A2(_09594_),
    .A3(_04700_),
    .B1(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__a31o_1 _28734_ (.A1(_04721_),
    .A2(_09594_),
    .A3(_04700_),
    .B1(_04824_),
    .X(_04826_));
 sky130_fd_sc_hd__a32oi_1 _28735_ (.A1(net171),
    .A2(_04722_),
    .A3(_04724_),
    .B1(_04729_),
    .B2(_04823_),
    .Y(_04827_));
 sky130_fd_sc_hd__a211oi_4 _28736_ (.A1(_04735_),
    .A2(_04729_),
    .B1(_04730_),
    .C1(_04825_),
    .Y(_04828_));
 sky130_fd_sc_hd__o211ai_4 _28737_ (.A1(_04736_),
    .A2(_04728_),
    .B1(_04731_),
    .C1(_04826_),
    .Y(_04829_));
 sky130_fd_sc_hd__and4_1 _28738_ (.A(_04822_),
    .B(_04616_),
    .C(_04612_),
    .D(_04332_),
    .X(_04830_));
 sky130_fd_sc_hd__nand3_1 _28739_ (.A(_04332_),
    .B(_04731_),
    .C(_04823_),
    .Y(_04831_));
 sky130_fd_sc_hd__nand3_4 _28740_ (.A(_04830_),
    .B(_04731_),
    .C(_04729_),
    .Y(_04834_));
 sky130_fd_sc_hd__inv_2 _28741_ (.A(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__a21oi_2 _28742_ (.A1(_04829_),
    .A2(_04834_),
    .B1(_04820_),
    .Y(_04836_));
 sky130_fd_sc_hd__o211ai_1 _28743_ (.A1(_04831_),
    .A2(_04728_),
    .B1(_04820_),
    .C1(_04829_),
    .Y(_04837_));
 sky130_fd_sc_hd__o21ai_2 _28744_ (.A1(net141),
    .A2(net139),
    .B1(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__a311o_2 _28745_ (.A1(net132),
    .A2(_04806_),
    .A3(_04807_),
    .B1(net130),
    .C1(_04797_),
    .X(_04839_));
 sky130_fd_sc_hd__a22oi_1 _28746_ (.A1(_04817_),
    .A2(_04819_),
    .B1(_04829_),
    .B2(_04834_),
    .Y(_04840_));
 sky130_fd_sc_hd__o22ai_2 _28747_ (.A1(_04816_),
    .A2(_04818_),
    .B1(_04828_),
    .B2(_04835_),
    .Y(_04841_));
 sky130_fd_sc_hd__o21ai_4 _28748_ (.A1(_10027_),
    .A2(_04814_),
    .B1(_04834_),
    .Y(_04842_));
 sky130_fd_sc_hd__o211ai_2 _28749_ (.A1(_04814_),
    .A2(_10027_),
    .B1(_04834_),
    .C1(_04829_),
    .Y(_04843_));
 sky130_fd_sc_hd__a211oi_1 _28750_ (.A1(_04740_),
    .A2(_04827_),
    .B1(_04816_),
    .C1(_04842_),
    .Y(_04845_));
 sky130_fd_sc_hd__o221ai_4 _28751_ (.A1(net141),
    .A2(net139),
    .B1(_04816_),
    .B2(_04843_),
    .C1(_04841_),
    .Y(_04846_));
 sky130_fd_sc_hd__o31a_2 _28752_ (.A1(_10479_),
    .A2(_04840_),
    .A3(_04845_),
    .B1(_04839_),
    .X(_04847_));
 sky130_fd_sc_hd__o221a_1 _28753_ (.A1(net130),
    .A2(_04814_),
    .B1(_04836_),
    .B2(_04838_),
    .C1(_10953_),
    .X(_04848_));
 sky130_fd_sc_hd__or3_1 _28754_ (.A(net137),
    .B(net134),
    .C(_04847_),
    .X(_04849_));
 sky130_fd_sc_hd__o311a_1 _28755_ (.A1(_10479_),
    .A2(_04840_),
    .A3(_04845_),
    .B1(_04839_),
    .C1(_09594_),
    .X(_04850_));
 sky130_fd_sc_hd__nand3_4 _28756_ (.A(_04846_),
    .B(_09594_),
    .C(_04839_),
    .Y(_04851_));
 sky130_fd_sc_hd__o221a_1 _28757_ (.A1(net130),
    .A2(_04814_),
    .B1(_04836_),
    .B2(_04838_),
    .C1(net171),
    .X(_04852_));
 sky130_fd_sc_hd__o221ai_4 _28758_ (.A1(net130),
    .A2(_04814_),
    .B1(_04836_),
    .B2(_04838_),
    .C1(net171),
    .Y(_04853_));
 sky130_fd_sc_hd__o211ai_2 _28759_ (.A1(_04624_),
    .A2(net176),
    .B1(_04751_),
    .C1(_04750_),
    .Y(_04854_));
 sky130_fd_sc_hd__o21ai_4 _28760_ (.A1(_09139_),
    .A2(_04743_),
    .B1(_04854_),
    .Y(_04856_));
 sky130_fd_sc_hd__a21oi_2 _28761_ (.A1(_04851_),
    .A2(_04853_),
    .B1(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__a21o_1 _28762_ (.A1(_04851_),
    .A2(_04853_),
    .B1(_04856_),
    .X(_04858_));
 sky130_fd_sc_hd__nand2_1 _28763_ (.A(_04853_),
    .B(_04856_),
    .Y(_04859_));
 sky130_fd_sc_hd__nand3_2 _28764_ (.A(_04851_),
    .B(_04853_),
    .C(_04856_),
    .Y(_04860_));
 sky130_fd_sc_hd__a31o_2 _28765_ (.A1(_04851_),
    .A2(_04853_),
    .A3(_04856_),
    .B1(_10953_),
    .X(_04861_));
 sky130_fd_sc_hd__o211ai_1 _28766_ (.A1(_04859_),
    .A2(_04850_),
    .B1(_10954_),
    .C1(_04858_),
    .Y(_04862_));
 sky130_fd_sc_hd__o22a_1 _28767_ (.A1(_10954_),
    .A2(_04847_),
    .B1(_04857_),
    .B2(_04861_),
    .X(_04863_));
 sky130_fd_sc_hd__o22ai_1 _28768_ (.A1(_10954_),
    .A2(_04847_),
    .B1(_04857_),
    .B2(_04861_),
    .Y(_04864_));
 sky130_fd_sc_hd__o221ai_4 _28769_ (.A1(_08313_),
    .A2(_04639_),
    .B1(_08730_),
    .B2(_04761_),
    .C1(_04655_),
    .Y(_04865_));
 sky130_fd_sc_hd__o21ai_1 _28770_ (.A1(_04857_),
    .A2(_04861_),
    .B1(_09139_),
    .Y(_04867_));
 sky130_fd_sc_hd__o221a_1 _28771_ (.A1(_10954_),
    .A2(_04847_),
    .B1(_04857_),
    .B2(_04861_),
    .C1(_09139_),
    .X(_04868_));
 sky130_fd_sc_hd__o221ai_4 _28772_ (.A1(_10954_),
    .A2(_04847_),
    .B1(_04857_),
    .B2(_04861_),
    .C1(_09139_),
    .Y(_04869_));
 sky130_fd_sc_hd__a2bb2oi_2 _28773_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_04849_),
    .B2(_04862_),
    .Y(_04870_));
 sky130_fd_sc_hd__o21ai_1 _28774_ (.A1(net194),
    .A2(net190),
    .B1(_04864_),
    .Y(_04871_));
 sky130_fd_sc_hd__o2111ai_1 _28775_ (.A1(net176),
    .A2(_04760_),
    .B1(_04865_),
    .C1(_04869_),
    .D1(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__o2bb2ai_1 _28776_ (.A1_N(_04763_),
    .A2_N(_04865_),
    .B1(_04868_),
    .B2(_04870_),
    .Y(_04873_));
 sky130_fd_sc_hd__o211ai_2 _28777_ (.A1(_11459_),
    .A2(net129),
    .B1(_04872_),
    .C1(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__o21ai_2 _28778_ (.A1(_11465_),
    .A2(_04863_),
    .B1(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__o21ai_2 _28779_ (.A1(_08724_),
    .A2(net196),
    .B1(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__inv_2 _28780_ (.A(_04876_),
    .Y(_04878_));
 sky130_fd_sc_hd__o211a_1 _28781_ (.A1(_11465_),
    .A2(_04863_),
    .B1(_08730_),
    .C1(_04874_),
    .X(_04879_));
 sky130_fd_sc_hd__o211ai_2 _28782_ (.A1(_04878_),
    .A2(_04879_),
    .B1(_04770_),
    .C1(_04780_),
    .Y(_04880_));
 sky130_fd_sc_hd__a21oi_1 _28783_ (.A1(_04880_),
    .A2(net133),
    .B1(_04875_),
    .Y(_04881_));
 sky130_fd_sc_hd__or3_1 _28784_ (.A(_05051_),
    .B(_04881_),
    .C(_04784_),
    .X(_04882_));
 sky130_fd_sc_hd__o21ai_1 _28785_ (.A1(_05051_),
    .A2(_04784_),
    .B1(_04881_),
    .Y(_04883_));
 sky130_fd_sc_hd__and2_1 _28786_ (.A(_04882_),
    .B(_04883_),
    .X(net116));
 sky130_fd_sc_hd__a2111o_1 _28787_ (.A1(net133),
    .A2(_04880_),
    .B1(_04875_),
    .C1(_04783_),
    .D1(_04665_),
    .X(_04884_));
 sky130_fd_sc_hd__o21ai_4 _28788_ (.A1(_10970_),
    .A2(_04785_),
    .B1(_11471_),
    .Y(_04885_));
 sky130_fd_sc_hd__o21ai_4 _28789_ (.A1(_04885_),
    .A2(_04792_),
    .B1(net144),
    .Y(_04886_));
 sky130_fd_sc_hd__or3_1 _28790_ (.A(net142),
    .B(_09573_),
    .C(_04886_),
    .X(_04888_));
 sky130_fd_sc_hd__o21ai_2 _28791_ (.A1(_10965_),
    .A2(_10967_),
    .B1(_04886_),
    .Y(_04889_));
 sky130_fd_sc_hd__o211ai_4 _28792_ (.A1(_04885_),
    .A2(_04792_),
    .B1(_10971_),
    .C1(net144),
    .Y(_04890_));
 sky130_fd_sc_hd__nand2_1 _28793_ (.A(_04889_),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__o211ai_2 _28794_ (.A1(net152),
    .A2(_04698_),
    .B1(_04719_),
    .C1(_04801_),
    .Y(_04892_));
 sky130_fd_sc_hd__o211ai_1 _28795_ (.A1(_04802_),
    .A2(_04805_),
    .B1(_04891_),
    .C1(_04801_),
    .Y(_04893_));
 sky130_fd_sc_hd__o2111ai_4 _28796_ (.A1(_10492_),
    .A2(_04796_),
    .B1(_04889_),
    .C1(_04890_),
    .D1(_04892_),
    .Y(_04894_));
 sky130_fd_sc_hd__nand3_2 _28797_ (.A(net132),
    .B(_04893_),
    .C(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__o21ai_2 _28798_ (.A1(net132),
    .A2(_04886_),
    .B1(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__inv_2 _28799_ (.A(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__a2bb2oi_1 _28800_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_04888_),
    .B2(_04895_),
    .Y(_04899_));
 sky130_fd_sc_hd__a2bb2o_1 _28801_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_04888_),
    .B2(_04895_),
    .X(_04900_));
 sky130_fd_sc_hd__o211a_1 _28802_ (.A1(net132),
    .A2(_04886_),
    .B1(_10491_),
    .C1(_04895_),
    .X(_04901_));
 sky130_fd_sc_hd__o211ai_2 _28803_ (.A1(net132),
    .A2(_04886_),
    .B1(_10491_),
    .C1(_04895_),
    .Y(_04902_));
 sky130_fd_sc_hd__nor2_1 _28804_ (.A(_04899_),
    .B(_04901_),
    .Y(_04903_));
 sky130_fd_sc_hd__o21ai_2 _28805_ (.A1(_04842_),
    .A2(_04828_),
    .B1(_04817_),
    .Y(_04904_));
 sky130_fd_sc_hd__o2111ai_1 _28806_ (.A1(_04842_),
    .A2(_04828_),
    .B1(_04817_),
    .C1(_04902_),
    .D1(_04900_),
    .Y(_04905_));
 sky130_fd_sc_hd__o21ai_1 _28807_ (.A1(_04899_),
    .A2(_04901_),
    .B1(_04904_),
    .Y(_04906_));
 sky130_fd_sc_hd__o211ai_1 _28808_ (.A1(net141),
    .A2(net139),
    .B1(_04905_),
    .C1(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__o221a_2 _28809_ (.A1(net152),
    .A2(_04815_),
    .B1(_04899_),
    .B2(_04901_),
    .C1(_04843_),
    .X(_04908_));
 sky130_fd_sc_hd__o2bb2ai_4 _28810_ (.A1_N(_04903_),
    .A2_N(_04904_),
    .B1(net141),
    .B2(net139),
    .Y(_04910_));
 sky130_fd_sc_hd__o22ai_4 _28811_ (.A1(net130),
    .A2(_04897_),
    .B1(_04908_),
    .B2(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__o22a_2 _28812_ (.A1(net130),
    .A2(_04897_),
    .B1(_04908_),
    .B2(_04910_),
    .X(_04912_));
 sky130_fd_sc_hd__o211a_1 _28813_ (.A1(net130),
    .A2(_04896_),
    .B1(_04907_),
    .C1(_10027_),
    .X(_04913_));
 sky130_fd_sc_hd__o21ai_4 _28814_ (.A1(net170),
    .A2(net168),
    .B1(_04911_),
    .Y(_04914_));
 sky130_fd_sc_hd__o221ai_4 _28815_ (.A1(net130),
    .A2(_04897_),
    .B1(_04908_),
    .B2(_04910_),
    .C1(net152),
    .Y(_04915_));
 sky130_fd_sc_hd__a21oi_1 _28816_ (.A1(_04624_),
    .A2(net176),
    .B1(_04482_),
    .Y(_04916_));
 sky130_fd_sc_hd__nor3_1 _28817_ (.A(_04628_),
    .B(_04482_),
    .C(_04626_),
    .Y(_04917_));
 sky130_fd_sc_hd__o2111a_1 _28818_ (.A1(net176),
    .A2(_04624_),
    .B1(_04916_),
    .C1(_04750_),
    .D1(_04747_),
    .X(_04918_));
 sky130_fd_sc_hd__nand3_2 _28819_ (.A(_04747_),
    .B(_04917_),
    .C(_04750_),
    .Y(_04919_));
 sky130_fd_sc_hd__a31oi_2 _28820_ (.A1(_04846_),
    .A2(_09594_),
    .A3(_04839_),
    .B1(_04919_),
    .Y(_04921_));
 sky130_fd_sc_hd__a21oi_1 _28821_ (.A1(_04851_),
    .A2(_04918_),
    .B1(_04852_),
    .Y(_04922_));
 sky130_fd_sc_hd__a211oi_4 _28822_ (.A1(_04856_),
    .A2(_04851_),
    .B1(_04852_),
    .C1(_04921_),
    .Y(_04923_));
 sky130_fd_sc_hd__o211ai_4 _28823_ (.A1(_04919_),
    .A2(_04850_),
    .B1(_04853_),
    .C1(_04860_),
    .Y(_04924_));
 sky130_fd_sc_hd__o2111a_1 _28824_ (.A1(_04726_),
    .A2(_04748_),
    .B1(_04494_),
    .C1(_04630_),
    .D1(_04747_),
    .X(_04925_));
 sky130_fd_sc_hd__nand3_4 _28825_ (.A(_04925_),
    .B(_04853_),
    .C(_04851_),
    .Y(_04926_));
 sky130_fd_sc_hd__a22oi_2 _28826_ (.A1(_04914_),
    .A2(_04915_),
    .B1(_04924_),
    .B2(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__a22o_1 _28827_ (.A1(_04914_),
    .A2(_04915_),
    .B1(_04924_),
    .B2(_04926_),
    .X(_04928_));
 sky130_fd_sc_hd__o21ai_4 _28828_ (.A1(_10027_),
    .A2(_04911_),
    .B1(_04926_),
    .Y(_04929_));
 sky130_fd_sc_hd__o211ai_4 _28829_ (.A1(_04911_),
    .A2(_10027_),
    .B1(_04926_),
    .C1(_04924_),
    .Y(_04930_));
 sky130_fd_sc_hd__a211oi_1 _28830_ (.A1(_04922_),
    .A2(_04860_),
    .B1(_04913_),
    .C1(_04929_),
    .Y(_04932_));
 sky130_fd_sc_hd__o221ai_4 _28831_ (.A1(net137),
    .A2(net134),
    .B1(_04913_),
    .B2(_04930_),
    .C1(_04928_),
    .Y(_04933_));
 sky130_fd_sc_hd__or3_2 _28832_ (.A(net137),
    .B(net134),
    .C(_04912_),
    .X(_04934_));
 sky130_fd_sc_hd__o31ai_2 _28833_ (.A1(_10953_),
    .A2(_04927_),
    .A3(_04932_),
    .B1(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__a211o_1 _28834_ (.A1(_04933_),
    .A2(_04934_),
    .B1(_11459_),
    .C1(net129),
    .X(_04936_));
 sky130_fd_sc_hd__o311a_2 _28835_ (.A1(_10953_),
    .A2(_04927_),
    .A3(_04932_),
    .B1(_04934_),
    .C1(_09594_),
    .X(_04937_));
 sky130_fd_sc_hd__nand3_1 _28836_ (.A(_04933_),
    .B(_04934_),
    .C(_09594_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21oi_1 _28837_ (.A1(_04933_),
    .A2(_04934_),
    .B1(_09594_),
    .Y(_04939_));
 sky130_fd_sc_hd__o21ai_2 _28838_ (.A1(net189),
    .A2(net186),
    .B1(_04935_),
    .Y(_04940_));
 sky130_fd_sc_hd__o221a_1 _28839_ (.A1(_04760_),
    .A2(net176),
    .B1(_09140_),
    .B2(_04864_),
    .C1(_04865_),
    .X(_04941_));
 sky130_fd_sc_hd__a31oi_4 _28840_ (.A1(_04763_),
    .A2(_04865_),
    .A3(_04869_),
    .B1(_04870_),
    .Y(_04944_));
 sky130_fd_sc_hd__o21a_1 _28841_ (.A1(_04937_),
    .A2(_04939_),
    .B1(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__o21ai_1 _28842_ (.A1(_04937_),
    .A2(_04939_),
    .B1(_04944_),
    .Y(_04946_));
 sky130_fd_sc_hd__o2bb2ai_1 _28843_ (.A1_N(net171),
    .A2_N(_04935_),
    .B1(_04941_),
    .B2(_04870_),
    .Y(_04947_));
 sky130_fd_sc_hd__o22ai_1 _28844_ (.A1(_11459_),
    .A2(net129),
    .B1(_04937_),
    .B2(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__o211ai_2 _28845_ (.A1(_04937_),
    .A2(_04947_),
    .B1(_04946_),
    .C1(_11465_),
    .Y(_04949_));
 sky130_fd_sc_hd__o21ai_2 _28846_ (.A1(_04945_),
    .A2(_04948_),
    .B1(_04936_),
    .Y(_04950_));
 sky130_fd_sc_hd__inv_2 _28847_ (.A(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__a21oi_1 _28848_ (.A1(_04936_),
    .A2(_04949_),
    .B1(_09139_),
    .Y(_04952_));
 sky130_fd_sc_hd__a2bb2o_1 _28849_ (.A1_N(net194),
    .A2_N(net190),
    .B1(_04936_),
    .B2(_04949_),
    .X(_04953_));
 sky130_fd_sc_hd__o211ai_2 _28850_ (.A1(_09136_),
    .A2(_09138_),
    .B1(_04936_),
    .C1(_04949_),
    .Y(_04955_));
 sky130_fd_sc_hd__a31oi_1 _28851_ (.A1(_04770_),
    .A2(_04780_),
    .A3(_04876_),
    .B1(_04879_),
    .Y(_04956_));
 sky130_fd_sc_hd__a21oi_1 _28852_ (.A1(_04953_),
    .A2(_04955_),
    .B1(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__o21ai_1 _28853_ (.A1(_11944_),
    .A2(_04957_),
    .B1(_04951_),
    .Y(_04958_));
 sky130_fd_sc_hd__a21oi_1 _28854_ (.A1(_05119_),
    .A2(_04884_),
    .B1(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__and3_1 _28855_ (.A(_05119_),
    .B(_04884_),
    .C(_04958_),
    .X(_04960_));
 sky130_fd_sc_hd__nor2_1 _28856_ (.A(_04959_),
    .B(_04960_),
    .Y(net117));
 sky130_fd_sc_hd__o2111ai_2 _28857_ (.A1(_11944_),
    .A2(_04957_),
    .B1(_04951_),
    .C1(_04881_),
    .D1(_04784_),
    .Y(_04961_));
 sky130_fd_sc_hd__o21ai_1 _28858_ (.A1(_04832_),
    .A2(_04942_),
    .B1(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__o32a_1 _28859_ (.A1(_03399_),
    .A2(net24),
    .A3(_10962_),
    .B1(_10970_),
    .B2(_04886_),
    .X(_04963_));
 sky130_fd_sc_hd__a21oi_4 _28860_ (.A1(_04894_),
    .A2(_04963_),
    .B1(_09578_),
    .Y(_04965_));
 sky130_fd_sc_hd__o21a_1 _28861_ (.A1(_10477_),
    .A2(_10478_),
    .B1(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__a311o_2 _28862_ (.A1(_11471_),
    .A2(_04890_),
    .A3(_04894_),
    .B1(_10970_),
    .C1(_09578_),
    .X(_04967_));
 sky130_fd_sc_hd__a21o_1 _28863_ (.A1(_10966_),
    .A2(_10968_),
    .B1(_04965_),
    .X(_04968_));
 sky130_fd_sc_hd__xor2_1 _28864_ (.A(_10971_),
    .B(_04965_),
    .X(_04969_));
 sky130_fd_sc_hd__o211ai_4 _28865_ (.A1(_04842_),
    .A2(_04828_),
    .B1(_04817_),
    .C1(_04900_),
    .Y(_04970_));
 sky130_fd_sc_hd__a22oi_4 _28866_ (.A1(_04967_),
    .A2(_04968_),
    .B1(_04970_),
    .B2(_04902_),
    .Y(_04971_));
 sky130_fd_sc_hd__o211a_1 _28867_ (.A1(_10492_),
    .A2(_04896_),
    .B1(_04969_),
    .C1(_04970_),
    .X(_04972_));
 sky130_fd_sc_hd__o211ai_2 _28868_ (.A1(_10492_),
    .A2(_04896_),
    .B1(_04969_),
    .C1(_04970_),
    .Y(_04973_));
 sky130_fd_sc_hd__o21ai_1 _28869_ (.A1(net141),
    .A2(net139),
    .B1(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__o22ai_2 _28870_ (.A1(net141),
    .A2(net139),
    .B1(_04971_),
    .B2(_04972_),
    .Y(_04976_));
 sky130_fd_sc_hd__o2bb2a_2 _28871_ (.A1_N(_10479_),
    .A2_N(_04965_),
    .B1(_04971_),
    .B2(_04974_),
    .X(_04977_));
 sky130_fd_sc_hd__a2bb2o_1 _28872_ (.A1_N(_04971_),
    .A2_N(_04974_),
    .B1(_10479_),
    .B2(_04965_),
    .X(_04978_));
 sky130_fd_sc_hd__or3_1 _28873_ (.A(net137),
    .B(net134),
    .C(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__o22ai_4 _28874_ (.A1(net152),
    .A2(_04912_),
    .B1(_04929_),
    .B2(_04923_),
    .Y(_04980_));
 sky130_fd_sc_hd__o21ai_2 _28875_ (.A1(_04971_),
    .A2(_04974_),
    .B1(_10491_),
    .Y(_04981_));
 sky130_fd_sc_hd__a21oi_1 _28876_ (.A1(_10479_),
    .A2(_04965_),
    .B1(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__o21ai_1 _28877_ (.A1(net164),
    .A2(_10490_),
    .B1(_04977_),
    .Y(_04983_));
 sky130_fd_sc_hd__o211a_1 _28878_ (.A1(_04965_),
    .A2(net130),
    .B1(_10492_),
    .C1(_04976_),
    .X(_04984_));
 sky130_fd_sc_hd__o211ai_2 _28879_ (.A1(_04965_),
    .A2(net130),
    .B1(_10492_),
    .C1(_04976_),
    .Y(_04985_));
 sky130_fd_sc_hd__o21ai_2 _28880_ (.A1(_04966_),
    .A2(_04981_),
    .B1(_04985_),
    .Y(_04987_));
 sky130_fd_sc_hd__o2111ai_1 _28881_ (.A1(_04929_),
    .A2(_04923_),
    .B1(_04914_),
    .C1(_04985_),
    .D1(_04983_),
    .Y(_04988_));
 sky130_fd_sc_hd__o21ai_1 _28882_ (.A1(_04982_),
    .A2(_04984_),
    .B1(_04980_),
    .Y(_04989_));
 sky130_fd_sc_hd__o211ai_2 _28883_ (.A1(net137),
    .A2(net134),
    .B1(_04988_),
    .C1(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__and3_1 _28884_ (.A(_10950_),
    .B(_10952_),
    .C(_04978_),
    .X(_04991_));
 sky130_fd_sc_hd__a21oi_4 _28885_ (.A1(_04914_),
    .A2(_04930_),
    .B1(_04987_),
    .Y(_04992_));
 sky130_fd_sc_hd__o221ai_4 _28886_ (.A1(net152),
    .A2(_04912_),
    .B1(_04929_),
    .B2(_04923_),
    .C1(_04987_),
    .Y(_04993_));
 sky130_fd_sc_hd__o21ai_4 _28887_ (.A1(net137),
    .A2(net134),
    .B1(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__o22ai_4 _28888_ (.A1(_10954_),
    .A2(_04977_),
    .B1(_04992_),
    .B2(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__inv_2 _28889_ (.A(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__and3_1 _28890_ (.A(_10027_),
    .B(_04979_),
    .C(_04990_),
    .X(_04998_));
 sky130_fd_sc_hd__o211ai_4 _28891_ (.A1(net170),
    .A2(net168),
    .B1(_04979_),
    .C1(_04990_),
    .Y(_04999_));
 sky130_fd_sc_hd__o22ai_1 _28892_ (.A1(net167),
    .A2(_10024_),
    .B1(_04992_),
    .B2(_04994_),
    .Y(_05000_));
 sky130_fd_sc_hd__o221ai_4 _28893_ (.A1(_10954_),
    .A2(_04977_),
    .B1(_04992_),
    .B2(_04994_),
    .C1(net152),
    .Y(_05001_));
 sky130_fd_sc_hd__o21a_1 _28894_ (.A1(_04991_),
    .A2(_05000_),
    .B1(_04999_),
    .X(_05002_));
 sky130_fd_sc_hd__o21ai_1 _28895_ (.A1(_04991_),
    .A2(_05000_),
    .B1(_04999_),
    .Y(_05003_));
 sky130_fd_sc_hd__o2111a_1 _28896_ (.A1(_04642_),
    .A2(_04638_),
    .B1(_04641_),
    .C1(_04763_),
    .D1(_04764_),
    .X(_05004_));
 sky130_fd_sc_hd__o211a_1 _28897_ (.A1(_04848_),
    .A2(_04867_),
    .B1(_05004_),
    .C1(_04871_),
    .X(_05005_));
 sky130_fd_sc_hd__nand2_1 _28898_ (.A(_04938_),
    .B(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__o211ai_4 _28899_ (.A1(_04944_),
    .A2(_04937_),
    .B1(_04940_),
    .C1(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__and4_1 _28900_ (.A(_05004_),
    .B(_04871_),
    .C(_04869_),
    .D(_04652_),
    .X(_05009_));
 sky130_fd_sc_hd__nand3_4 _28901_ (.A(_04938_),
    .B(_04940_),
    .C(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__a21oi_1 _28902_ (.A1(_05007_),
    .A2(_05010_),
    .B1(_05003_),
    .Y(_05011_));
 sky130_fd_sc_hd__a31o_1 _28903_ (.A1(_05003_),
    .A2(_05007_),
    .A3(_05010_),
    .B1(_11464_),
    .X(_05012_));
 sky130_fd_sc_hd__or3_1 _28904_ (.A(_11459_),
    .B(net129),
    .C(_04996_),
    .X(_05013_));
 sky130_fd_sc_hd__a22oi_2 _28905_ (.A1(_04999_),
    .A2(_05001_),
    .B1(_05007_),
    .B2(_05010_),
    .Y(_05014_));
 sky130_fd_sc_hd__a21o_1 _28906_ (.A1(_05007_),
    .A2(_05010_),
    .B1(_05002_),
    .X(_05015_));
 sky130_fd_sc_hd__o211ai_2 _28907_ (.A1(_04995_),
    .A2(_10027_),
    .B1(_05010_),
    .C1(_05007_),
    .Y(_05016_));
 sky130_fd_sc_hd__o2111a_1 _28908_ (.A1(_10027_),
    .A2(_04995_),
    .B1(_04999_),
    .C1(_05007_),
    .D1(_05010_),
    .X(_05017_));
 sky130_fd_sc_hd__o221ai_1 _28909_ (.A1(_11459_),
    .A2(net129),
    .B1(_04998_),
    .B2(_05016_),
    .C1(_05015_),
    .Y(_05018_));
 sky130_fd_sc_hd__o31a_1 _28910_ (.A1(_11464_),
    .A2(_05014_),
    .A3(_05017_),
    .B1(_05013_),
    .X(_05020_));
 sky130_fd_sc_hd__o311a_1 _28911_ (.A1(_11464_),
    .A2(_05014_),
    .A3(_05017_),
    .B1(_05013_),
    .C1(_09594_),
    .X(_05021_));
 sky130_fd_sc_hd__nand3_1 _28912_ (.A(_05018_),
    .B(_09594_),
    .C(_05013_),
    .Y(_05022_));
 sky130_fd_sc_hd__o221ai_4 _28913_ (.A1(_11465_),
    .A2(_04995_),
    .B1(_05011_),
    .B2(_05012_),
    .C1(net171),
    .Y(_05023_));
 sky130_fd_sc_hd__nand2_1 _28914_ (.A(_05022_),
    .B(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__a21oi_1 _28915_ (.A1(_04956_),
    .A2(_04955_),
    .B1(_04952_),
    .Y(_05025_));
 sky130_fd_sc_hd__a21boi_1 _28916_ (.A1(_05022_),
    .A2(_05023_),
    .B1_N(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__o21ai_2 _28917_ (.A1(_11944_),
    .A2(_05026_),
    .B1(_05020_),
    .Y(_05027_));
 sky130_fd_sc_hd__xnor2_1 _28918_ (.A(_04962_),
    .B(_05027_),
    .Y(net118));
 sky130_fd_sc_hd__nor2_1 _28919_ (.A(_04961_),
    .B(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__o22a_1 _28920_ (.A1(_04832_),
    .A2(_04942_),
    .B1(_04961_),
    .B2(_05027_),
    .X(_05030_));
 sky130_fd_sc_hd__a31oi_2 _28921_ (.A1(_11471_),
    .A2(_04967_),
    .A3(_04973_),
    .B1(_10479_),
    .Y(_05031_));
 sky130_fd_sc_hd__a311o_2 _28922_ (.A1(_11471_),
    .A2(_04967_),
    .A3(_04973_),
    .B1(_10954_),
    .C1(_10479_),
    .X(_05032_));
 sky130_fd_sc_hd__xor2_1 _28923_ (.A(_10971_),
    .B(_05031_),
    .X(_05033_));
 sky130_fd_sc_hd__xor2_1 _28924_ (.A(_10970_),
    .B(_05031_),
    .X(_05034_));
 sky130_fd_sc_hd__o21ai_1 _28925_ (.A1(_10492_),
    .A2(_04978_),
    .B1(_04980_),
    .Y(_05035_));
 sky130_fd_sc_hd__o221ai_4 _28926_ (.A1(_04966_),
    .A2(_04981_),
    .B1(_04984_),
    .B2(_04980_),
    .C1(_05033_),
    .Y(_05036_));
 sky130_fd_sc_hd__o211ai_2 _28927_ (.A1(_10491_),
    .A2(_04977_),
    .B1(_05034_),
    .C1(_05035_),
    .Y(_05037_));
 sky130_fd_sc_hd__o211ai_4 _28928_ (.A1(net137),
    .A2(net134),
    .B1(_05036_),
    .C1(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__a21oi_4 _28929_ (.A1(_05032_),
    .A2(_05038_),
    .B1(_11465_),
    .Y(_05039_));
 sky130_fd_sc_hd__a2bb2oi_2 _28930_ (.A1_N(_10487_),
    .A2_N(net165),
    .B1(_05032_),
    .B2(_05038_),
    .Y(_05041_));
 sky130_fd_sc_hd__a211o_1 _28931_ (.A1(_05032_),
    .A2(_05038_),
    .B1(net164),
    .C1(_10490_),
    .X(_05042_));
 sky130_fd_sc_hd__a31oi_1 _28932_ (.A1(_10954_),
    .A2(_05036_),
    .A3(_05037_),
    .B1(_10492_),
    .Y(_05043_));
 sky130_fd_sc_hd__and3_1 _28933_ (.A(_05038_),
    .B(_10491_),
    .C(_05032_),
    .X(_05044_));
 sky130_fd_sc_hd__a21oi_1 _28934_ (.A1(_05032_),
    .A2(_05043_),
    .B1(_05041_),
    .Y(_05045_));
 sky130_fd_sc_hd__o2bb2ai_1 _28935_ (.A1_N(_05007_),
    .A2_N(_05010_),
    .B1(net152),
    .B2(_04996_),
    .Y(_05046_));
 sky130_fd_sc_hd__a31oi_1 _28936_ (.A1(_05001_),
    .A2(_05007_),
    .A3(_05010_),
    .B1(_04998_),
    .Y(_05047_));
 sky130_fd_sc_hd__o211ai_4 _28937_ (.A1(_10027_),
    .A2(_04995_),
    .B1(_05045_),
    .C1(_05046_),
    .Y(_05048_));
 sky130_fd_sc_hd__o221ai_4 _28938_ (.A1(net152),
    .A2(_04996_),
    .B1(_05041_),
    .B2(_05044_),
    .C1(_05016_),
    .Y(_05049_));
 sky130_fd_sc_hd__o311a_1 _28939_ (.A1(_05041_),
    .A2(_05044_),
    .A3(_05047_),
    .B1(_05049_),
    .C1(_11465_),
    .X(_05050_));
 sky130_fd_sc_hd__a31oi_4 _28940_ (.A1(_11465_),
    .A2(_05048_),
    .A3(_05049_),
    .B1(_05039_),
    .Y(_05053_));
 sky130_fd_sc_hd__o21ai_4 _28941_ (.A1(_05039_),
    .A2(_05050_),
    .B1(_10027_),
    .Y(_05054_));
 sky130_fd_sc_hd__a311o_1 _28942_ (.A1(_11465_),
    .A2(_05048_),
    .A3(_05049_),
    .B1(_05039_),
    .C1(_10027_),
    .X(_05055_));
 sky130_fd_sc_hd__nor3b_1 _28943_ (.A(_04879_),
    .B(_04772_),
    .C_N(_04876_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand3b_1 _28944_ (.A_N(_04879_),
    .B(_04771_),
    .C(_04876_),
    .Y(_05057_));
 sky130_fd_sc_hd__a21oi_1 _28945_ (.A1(_09140_),
    .A2(_04950_),
    .B1(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__nand3_1 _28946_ (.A(_04953_),
    .B(_05056_),
    .C(_04955_),
    .Y(_05059_));
 sky130_fd_sc_hd__o211ai_1 _28947_ (.A1(_09140_),
    .A2(_04950_),
    .B1(_05058_),
    .C1(_05022_),
    .Y(_05060_));
 sky130_fd_sc_hd__o211a_2 _28948_ (.A1(_05025_),
    .A2(_05021_),
    .B1(_05023_),
    .C1(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__o211ai_1 _28949_ (.A1(_05025_),
    .A2(_05021_),
    .B1(_05023_),
    .C1(_05060_),
    .Y(_05062_));
 sky130_fd_sc_hd__nand4_2 _28950_ (.A(_04953_),
    .B(_05056_),
    .C(_04955_),
    .D(_04779_),
    .Y(_05064_));
 sky130_fd_sc_hd__nand4b_1 _28951_ (.A_N(_05059_),
    .B(_05023_),
    .C(_05022_),
    .D(_04779_),
    .Y(_05065_));
 sky130_fd_sc_hd__o211ai_2 _28952_ (.A1(_05024_),
    .A2(_05064_),
    .B1(_05055_),
    .C1(_05054_),
    .Y(_05066_));
 sky130_fd_sc_hd__a22o_1 _28953_ (.A1(_05054_),
    .A2(_05055_),
    .B1(_05062_),
    .B2(_05065_),
    .X(_05067_));
 sky130_fd_sc_hd__o211ai_4 _28954_ (.A1(_05061_),
    .A2(_05066_),
    .B1(net133),
    .C1(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__o211a_1 _28955_ (.A1(_05051_),
    .A2(_05028_),
    .B1(_05053_),
    .C1(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__a211oi_1 _28956_ (.A1(_05068_),
    .A2(_05053_),
    .B1(_05028_),
    .C1(_05051_),
    .Y(_05070_));
 sky130_fd_sc_hd__nor2_1 _28957_ (.A(_05069_),
    .B(_05070_),
    .Y(net119));
 sky130_fd_sc_hd__o2bb2a_1 _28958_ (.A1_N(_05031_),
    .A2_N(_10971_),
    .B1(net24),
    .B2(_11469_),
    .X(_05071_));
 sky130_fd_sc_hd__a21oi_4 _28959_ (.A1(_05036_),
    .A2(_05071_),
    .B1(_10953_),
    .Y(_05072_));
 sky130_fd_sc_hd__and3_1 _28960_ (.A(_05072_),
    .B(_10968_),
    .C(_10966_),
    .X(_05074_));
 sky130_fd_sc_hd__xor2_2 _28961_ (.A(_10970_),
    .B(_05072_),
    .X(_05075_));
 sky130_fd_sc_hd__inv_2 _28962_ (.A(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__o21ai_1 _28963_ (.A1(_05044_),
    .A2(_05047_),
    .B1(_05042_),
    .Y(_05077_));
 sky130_fd_sc_hd__a21oi_2 _28964_ (.A1(_05042_),
    .A2(_05048_),
    .B1(_05075_),
    .Y(_05078_));
 sky130_fd_sc_hd__nand2_1 _28965_ (.A(_05077_),
    .B(_05076_),
    .Y(_05079_));
 sky130_fd_sc_hd__a31oi_2 _28966_ (.A1(_05042_),
    .A2(_05048_),
    .A3(_05075_),
    .B1(_11464_),
    .Y(_05080_));
 sky130_fd_sc_hd__a22oi_2 _28967_ (.A1(_11464_),
    .A2(_05072_),
    .B1(_05080_),
    .B2(_05079_),
    .Y(_05081_));
 sky130_fd_sc_hd__a22o_1 _28968_ (.A1(_11464_),
    .A2(_05072_),
    .B1(_05080_),
    .B2(_05079_),
    .X(_05082_));
 sky130_fd_sc_hd__nor2_1 _28969_ (.A(net133),
    .B(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__o2bb2ai_2 _28970_ (.A1_N(net152),
    .A2_N(_05053_),
    .B1(_05064_),
    .B2(_05024_),
    .Y(_05085_));
 sky130_fd_sc_hd__o22ai_1 _28971_ (.A1(net152),
    .A2(_05053_),
    .B1(_05085_),
    .B2(_05061_),
    .Y(_05086_));
 sky130_fd_sc_hd__o21ai_2 _28972_ (.A1(net164),
    .A2(_10490_),
    .B1(_05081_),
    .Y(_05087_));
 sky130_fd_sc_hd__o21ai_1 _28973_ (.A1(_10487_),
    .A2(net165),
    .B1(_05082_),
    .Y(_05088_));
 sky130_fd_sc_hd__o2111ai_2 _28974_ (.A1(_05085_),
    .A2(_05061_),
    .B1(_05054_),
    .C1(_05088_),
    .D1(_05087_),
    .Y(_05089_));
 sky130_fd_sc_hd__nand3_1 _28975_ (.A(_05086_),
    .B(_05087_),
    .C(_05088_),
    .Y(_05090_));
 sky130_fd_sc_hd__a21oi_1 _28976_ (.A1(_05089_),
    .A2(net133),
    .B1(_05083_),
    .Y(_05091_));
 sky130_fd_sc_hd__a21oi_1 _28977_ (.A1(_05068_),
    .A2(_05053_),
    .B1(_05051_),
    .Y(_05092_));
 sky130_fd_sc_hd__a31o_1 _28978_ (.A1(_05068_),
    .A2(_05053_),
    .A3(_05028_),
    .B1(_05051_),
    .X(_05093_));
 sky130_fd_sc_hd__a31oi_2 _28979_ (.A1(_05068_),
    .A2(_05053_),
    .A3(_05028_),
    .B1(_05051_),
    .Y(_05094_));
 sky130_fd_sc_hd__xor2_1 _28980_ (.A(_05091_),
    .B(_05094_),
    .X(net121));
 sky130_fd_sc_hd__o21a_1 _28981_ (.A1(_04832_),
    .A2(_04942_),
    .B1(_05091_),
    .X(_05096_));
 sky130_fd_sc_hd__a211o_1 _28982_ (.A1(_05089_),
    .A2(net133),
    .B1(_05051_),
    .C1(_05083_),
    .X(_05097_));
 sky130_fd_sc_hd__a21oi_1 _28983_ (.A1(_05119_),
    .A2(_05091_),
    .B1(_05094_),
    .Y(_05098_));
 sky130_fd_sc_hd__a211oi_1 _28984_ (.A1(_05077_),
    .A2(_05076_),
    .B1(_05074_),
    .C1(_11470_),
    .Y(_05099_));
 sky130_fd_sc_hd__o32a_1 _28985_ (.A1(_11470_),
    .A2(_05074_),
    .A3(_05078_),
    .B1(net129),
    .B2(_11459_),
    .X(_05100_));
 sky130_fd_sc_hd__o21ai_1 _28986_ (.A1(_11464_),
    .A2(_05099_),
    .B1(_10970_),
    .Y(_05101_));
 sky130_fd_sc_hd__o311ai_4 _28987_ (.A1(_11470_),
    .A2(_05074_),
    .A3(_05078_),
    .B1(_11465_),
    .C1(_10971_),
    .Y(_05102_));
 sky130_fd_sc_hd__o221ai_2 _28988_ (.A1(_10491_),
    .A2(_05081_),
    .B1(_05085_),
    .B2(_05061_),
    .C1(_05054_),
    .Y(_05103_));
 sky130_fd_sc_hd__a22oi_1 _28989_ (.A1(_10492_),
    .A2(_05082_),
    .B1(_05101_),
    .B2(_05102_),
    .Y(_05104_));
 sky130_fd_sc_hd__a22oi_1 _28990_ (.A1(_05101_),
    .A2(_05102_),
    .B1(_05103_),
    .B2(_05087_),
    .Y(_05106_));
 sky130_fd_sc_hd__a21oi_1 _28991_ (.A1(_05090_),
    .A2(_05104_),
    .B1(_11944_),
    .Y(_05107_));
 sky130_fd_sc_hd__o22a_1 _28992_ (.A1(_11464_),
    .A2(_05099_),
    .B1(_11944_),
    .B2(_05106_),
    .X(_05108_));
 sky130_fd_sc_hd__a211o_1 _28993_ (.A1(_05097_),
    .A2(_05093_),
    .B1(_05107_),
    .C1(_05100_),
    .X(_05109_));
 sky130_fd_sc_hd__o41ai_1 _28994_ (.A1(_05030_),
    .A2(_05092_),
    .A3(_05096_),
    .A4(_05108_),
    .B1(_05109_),
    .Y(net122));
 sky130_fd_sc_hd__o22ai_1 _28995_ (.A1(_04832_),
    .A2(_04942_),
    .B1(_05100_),
    .B2(_05107_),
    .Y(_05110_));
 sky130_fd_sc_hd__o221ai_1 _28996_ (.A1(_10492_),
    .A2(_05082_),
    .B1(_05100_),
    .B2(_10971_),
    .C1(_05103_),
    .Y(_05111_));
 sky130_fd_sc_hd__a31o_1 _28997_ (.A1(_11471_),
    .A2(_05102_),
    .A3(_05111_),
    .B1(_11944_),
    .X(_05112_));
 sky130_fd_sc_hd__a31oi_1 _28998_ (.A1(_05110_),
    .A2(_05093_),
    .A3(_05097_),
    .B1(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__o211a_1 _28999_ (.A1(_05051_),
    .A2(_05108_),
    .B1(_05112_),
    .C1(_05098_),
    .X(_05114_));
 sky130_fd_sc_hd__nor2_1 _29000_ (.A(_05113_),
    .B(_05114_),
    .Y(net123));
 sky130_fd_sc_hd__nor2_1 _29001_ (.A(_05051_),
    .B(_05114_),
    .Y(net124));
 sky130_fd_sc_hd__clkbuf_16 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_8 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_8 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_8 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_16 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_8 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_6 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_6 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_8 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_8 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_12 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_8 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_6 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_8 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_6 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_6 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_6 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_16 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_8 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_4 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_8 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_8 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_6 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_4 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_6 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_4 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_4 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_2 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 output65 (.A(net65),
    .X(Product[0]));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(Product[10]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(Product[11]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(Product[12]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(Product[13]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(Product[14]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(Product[15]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(Product[16]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(Product[17]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(Product[18]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(Product[19]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(Product[1]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(Product[20]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(Product[21]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(Product[22]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(Product[23]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(Product[24]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(Product[25]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(Product[26]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(Product[27]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(Product[28]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(Product[29]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(Product[2]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(Product[30]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(Product[31]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(Product[32]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(Product[33]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(Product[34]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(Product[35]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(Product[36]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(Product[37]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(Product[38]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(Product[39]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(Product[3]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(Product[40]));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(Product[41]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(Product[42]));
 sky130_fd_sc_hd__buf_1 output102 (.A(net102),
    .X(Product[43]));
 sky130_fd_sc_hd__buf_1 output103 (.A(net103),
    .X(Product[44]));
 sky130_fd_sc_hd__buf_1 output104 (.A(net104),
    .X(Product[45]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(Product[46]));
 sky130_fd_sc_hd__buf_1 output106 (.A(net106),
    .X(Product[47]));
 sky130_fd_sc_hd__buf_1 output107 (.A(net107),
    .X(Product[48]));
 sky130_fd_sc_hd__buf_1 output108 (.A(net108),
    .X(Product[49]));
 sky130_fd_sc_hd__buf_1 output109 (.A(net109),
    .X(Product[4]));
 sky130_fd_sc_hd__buf_1 output110 (.A(net110),
    .X(Product[50]));
 sky130_fd_sc_hd__buf_1 output111 (.A(net111),
    .X(Product[51]));
 sky130_fd_sc_hd__buf_1 output112 (.A(net112),
    .X(Product[52]));
 sky130_fd_sc_hd__buf_1 output113 (.A(net113),
    .X(Product[53]));
 sky130_fd_sc_hd__buf_1 output114 (.A(net114),
    .X(Product[54]));
 sky130_fd_sc_hd__buf_1 output115 (.A(net115),
    .X(Product[55]));
 sky130_fd_sc_hd__buf_1 output116 (.A(net116),
    .X(Product[56]));
 sky130_fd_sc_hd__buf_1 output117 (.A(net117),
    .X(Product[57]));
 sky130_fd_sc_hd__buf_1 output118 (.A(net118),
    .X(Product[58]));
 sky130_fd_sc_hd__buf_1 output119 (.A(net119),
    .X(Product[59]));
 sky130_fd_sc_hd__buf_1 output120 (.A(net120),
    .X(Product[5]));
 sky130_fd_sc_hd__buf_1 output121 (.A(net121),
    .X(Product[60]));
 sky130_fd_sc_hd__buf_1 output122 (.A(net122),
    .X(Product[61]));
 sky130_fd_sc_hd__buf_1 output123 (.A(net123),
    .X(Product[62]));
 sky130_fd_sc_hd__buf_1 output124 (.A(net124),
    .X(Product[63]));
 sky130_fd_sc_hd__buf_1 output125 (.A(net125),
    .X(Product[6]));
 sky130_fd_sc_hd__buf_1 output126 (.A(net126),
    .X(Product[7]));
 sky130_fd_sc_hd__buf_1 output127 (.A(net127),
    .X(Product[8]));
 sky130_fd_sc_hd__buf_1 output128 (.A(net128),
    .X(Product[9]));
 sky130_fd_sc_hd__buf_12 max_cap129 (.A(_11461_),
    .X(net129));
 sky130_fd_sc_hd__buf_12 max_cap130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__buf_12 wire131 (.A(_10480_),
    .X(net131));
 sky130_fd_sc_hd__buf_12 max_cap132 (.A(_09579_),
    .X(net132));
 sky130_fd_sc_hd__buf_4 max_cap133 (.A(_11943_),
    .X(net133));
 sky130_fd_sc_hd__buf_8 max_cap134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_8 max_cap135 (.A(_10951_),
    .X(net135));
 sky130_fd_sc_hd__buf_8 max_cap136 (.A(_10951_),
    .X(net136));
 sky130_fd_sc_hd__buf_12 max_cap137 (.A(_10949_),
    .X(net137));
 sky130_fd_sc_hd__buf_8 max_cap138 (.A(_10475_),
    .X(net138));
 sky130_fd_sc_hd__buf_8 max_cap139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_8 max_cap140 (.A(_10475_),
    .X(net140));
 sky130_fd_sc_hd__buf_12 max_cap141 (.A(_10474_),
    .X(net141));
 sky130_fd_sc_hd__buf_12 max_cap142 (.A(_09571_),
    .X(net142));
 sky130_fd_sc_hd__buf_12 max_cap143 (.A(_09563_),
    .X(net143));
 sky130_fd_sc_hd__buf_12 max_cap144 (.A(_09563_),
    .X(net144));
 sky130_fd_sc_hd__buf_12 max_cap145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_12 max_cap146 (.A(_09125_),
    .X(net146));
 sky130_fd_sc_hd__buf_12 max_cap147 (.A(_09121_),
    .X(net147));
 sky130_fd_sc_hd__buf_12 max_cap148 (.A(_09120_),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_16 max_cap149 (.A(_08714_),
    .X(net149));
 sky130_fd_sc_hd__buf_12 max_cap150 (.A(_10491_),
    .X(net150));
 sky130_fd_sc_hd__buf_12 max_cap151 (.A(_10027_),
    .X(net151));
 sky130_fd_sc_hd__buf_12 wire152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__buf_12 max_cap153 (.A(_10026_),
    .X(net153));
 sky130_fd_sc_hd__buf_8 max_cap154 (.A(_09556_),
    .X(net154));
 sky130_fd_sc_hd__buf_8 max_cap155 (.A(_09556_),
    .X(net155));
 sky130_fd_sc_hd__buf_12 max_cap156 (.A(_09553_),
    .X(net156));
 sky130_fd_sc_hd__buf_8 max_cap157 (.A(_08709_),
    .X(net157));
 sky130_fd_sc_hd__buf_8 max_cap158 (.A(_08709_),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_16 max_cap159 (.A(_08300_),
    .X(net159));
 sky130_fd_sc_hd__buf_12 max_cap160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_12 max_cap161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__buf_12 max_cap162 (.A(_07916_),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_16 max_cap163 (.A(_07548_),
    .X(net163));
 sky130_fd_sc_hd__buf_12 max_cap164 (.A(_10489_),
    .X(net164));
 sky130_fd_sc_hd__buf_8 max_cap165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_8 max_cap166 (.A(_10488_),
    .X(net166));
 sky130_fd_sc_hd__buf_8 max_cap167 (.A(_10023_),
    .X(net167));
 sky130_fd_sc_hd__buf_8 max_cap168 (.A(_10022_),
    .X(net168));
 sky130_fd_sc_hd__buf_12 max_cap169 (.A(_10022_),
    .X(net169));
 sky130_fd_sc_hd__buf_12 max_cap170 (.A(_10021_),
    .X(net170));
 sky130_fd_sc_hd__buf_12 wire171 (.A(_09595_),
    .X(net171));
 sky130_fd_sc_hd__buf_12 max_cap172 (.A(_09594_),
    .X(net172));
 sky130_fd_sc_hd__buf_12 max_cap173 (.A(_09140_),
    .X(net173));
 sky130_fd_sc_hd__buf_12 max_cap174 (.A(_09139_),
    .X(net174));
 sky130_fd_sc_hd__buf_12 max_cap175 (.A(_08731_),
    .X(net175));
 sky130_fd_sc_hd__buf_12 max_cap176 (.A(_08731_),
    .X(net176));
 sky130_fd_sc_hd__buf_12 max_cap177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_12 max_cap178 (.A(_08730_),
    .X(net178));
 sky130_fd_sc_hd__buf_12 max_cap179 (.A(_08298_),
    .X(net179));
 sky130_fd_sc_hd__buf_8 max_cap180 (.A(_08296_),
    .X(net180));
 sky130_fd_sc_hd__buf_8 max_cap181 (.A(_08296_),
    .X(net181));
 sky130_fd_sc_hd__buf_12 max_cap182 (.A(_07914_),
    .X(net182));
 sky130_fd_sc_hd__buf_12 max_cap183 (.A(_07912_),
    .X(net183));
 sky130_fd_sc_hd__buf_12 max_cap184 (.A(_07546_),
    .X(net184));
 sky130_fd_sc_hd__buf_12 max_cap185 (.A(_07233_),
    .X(net185));
 sky130_fd_sc_hd__buf_8 max_cap186 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__buf_8 max_cap187 (.A(_09590_),
    .X(net187));
 sky130_fd_sc_hd__buf_8 max_cap188 (.A(_09590_),
    .X(net188));
 sky130_fd_sc_hd__buf_12 max_cap189 (.A(_09588_),
    .X(net189));
 sky130_fd_sc_hd__buf_8 max_cap190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_8 max_cap191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_6 max_cap192 (.A(_09135_),
    .X(net192));
 sky130_fd_sc_hd__buf_12 max_cap193 (.A(_09135_),
    .X(net193));
 sky130_fd_sc_hd__buf_12 max_cap194 (.A(_09134_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 max_cap195 (.A(_08729_),
    .X(net195));
 sky130_fd_sc_hd__buf_12 max_cap196 (.A(_08726_),
    .X(net196));
 sky130_fd_sc_hd__buf_12 max_cap197 (.A(_08314_),
    .X(net197));
 sky130_fd_sc_hd__buf_12 max_cap198 (.A(_08314_),
    .X(net198));
 sky130_fd_sc_hd__buf_12 max_cap199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_12 max_cap200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_12 max_cap201 (.A(_08313_),
    .X(net201));
 sky130_fd_sc_hd__buf_12 max_cap202 (.A(_07565_),
    .X(net202));
 sky130_fd_sc_hd__buf_8 max_cap203 (.A(_07229_),
    .X(net203));
 sky130_fd_sc_hd__buf_8 max_cap204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_8 max_cap205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__buf_12 max_cap206 (.A(_07229_),
    .X(net206));
 sky130_fd_sc_hd__buf_12 max_cap207 (.A(_07227_),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_16 wire208 (.A(_06903_),
    .X(net208));
 sky130_fd_sc_hd__buf_12 max_cap209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_12 max_cap210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_12 max_cap211 (.A(_06612_),
    .X(net211));
 sky130_fd_sc_hd__buf_12 max_cap212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__buf_12 max_cap213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__buf_12 max_cap214 (.A(_06293_),
    .X(net214));
 sky130_fd_sc_hd__buf_8 max_cap215 (.A(_08312_),
    .X(net215));
 sky130_fd_sc_hd__buf_12 max_cap216 (.A(_08309_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_8 max_cap217 (.A(_07562_),
    .X(net217));
 sky130_fd_sc_hd__buf_8 max_cap218 (.A(_07557_),
    .X(net218));
 sky130_fd_sc_hd__buf_8 max_cap219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__buf_8 wire220 (.A(_07557_),
    .X(net220));
 sky130_fd_sc_hd__buf_12 max_cap221 (.A(_07555_),
    .X(net221));
 sky130_fd_sc_hd__buf_12 max_cap222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_12 max_cap223 (.A(_07247_),
    .X(net223));
 sky130_fd_sc_hd__buf_12 max_cap224 (.A(_07246_),
    .X(net224));
 sky130_fd_sc_hd__buf_12 max_cap225 (.A(_06924_),
    .X(net225));
 sky130_fd_sc_hd__buf_12 max_cap226 (.A(_06924_),
    .X(net226));
 sky130_fd_sc_hd__buf_12 max_cap227 (.A(_06922_),
    .X(net227));
 sky130_fd_sc_hd__buf_12 max_cap228 (.A(_06901_),
    .X(net228));
 sky130_fd_sc_hd__buf_8 max_cap229 (.A(net231),
    .X(net229));
 sky130_fd_sc_hd__buf_8 max_cap230 (.A(_06899_),
    .X(net230));
 sky130_fd_sc_hd__buf_8 max_cap231 (.A(_06899_),
    .X(net231));
 sky130_fd_sc_hd__buf_12 max_cap232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_12 max_cap233 (.A(_06630_),
    .X(net233));
 sky130_fd_sc_hd__buf_12 max_cap234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__buf_12 max_cap235 (.A(_06629_),
    .X(net235));
 sky130_fd_sc_hd__buf_8 max_cap236 (.A(_06610_),
    .X(net236));
 sky130_fd_sc_hd__buf_8 max_cap237 (.A(_06610_),
    .X(net237));
 sky130_fd_sc_hd__buf_12 max_cap238 (.A(_06608_),
    .X(net238));
 sky130_fd_sc_hd__buf_8 max_cap239 (.A(_06291_),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_16 max_cap240 (.A(_05996_),
    .X(net240));
 sky130_fd_sc_hd__buf_12 wire241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_12 max_cap242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__buf_12 max_cap243 (.A(_05752_),
    .X(net243));
 sky130_fd_sc_hd__buf_12 max_cap244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__buf_12 max_cap245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_12 max_cap246 (.A(_05485_),
    .X(net246));
 sky130_fd_sc_hd__buf_6 max_cap247 (.A(_07245_),
    .X(net247));
 sky130_fd_sc_hd__buf_12 max_cap248 (.A(_07243_),
    .X(net248));
 sky130_fd_sc_hd__buf_8 max_cap249 (.A(_06920_),
    .X(net249));
 sky130_fd_sc_hd__buf_12 max_cap250 (.A(_06916_),
    .X(net250));
 sky130_fd_sc_hd__buf_12 max_cap251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_12 max_cap252 (.A(_06315_),
    .X(net252));
 sky130_fd_sc_hd__buf_12 max_cap253 (.A(_06014_),
    .X(net253));
 sky130_fd_sc_hd__buf_12 max_cap254 (.A(_06013_),
    .X(net254));
 sky130_fd_sc_hd__buf_8 wire255 (.A(net258),
    .X(net255));
 sky130_fd_sc_hd__buf_8 max_cap256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_8 max_cap257 (.A(_05992_),
    .X(net257));
 sky130_fd_sc_hd__buf_12 max_cap258 (.A(_05992_),
    .X(net258));
 sky130_fd_sc_hd__buf_12 max_cap259 (.A(_05990_),
    .X(net259));
 sky130_fd_sc_hd__buf_12 max_cap260 (.A(_05990_),
    .X(net260));
 sky130_fd_sc_hd__buf_12 max_cap261 (.A(_05768_),
    .X(net261));
 sky130_fd_sc_hd__buf_12 max_cap262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__buf_12 max_cap263 (.A(_05767_),
    .X(net263));
 sky130_fd_sc_hd__buf_12 max_cap264 (.A(_05751_),
    .X(net264));
 sky130_fd_sc_hd__buf_8 max_cap265 (.A(_05750_),
    .X(net265));
 sky130_fd_sc_hd__buf_12 max_cap266 (.A(_05750_),
    .X(net266));
 sky130_fd_sc_hd__buf_12 max_cap267 (.A(_05507_),
    .X(net267));
 sky130_fd_sc_hd__buf_8 max_cap268 (.A(_05483_),
    .X(net268));
 sky130_fd_sc_hd__buf_8 max_cap269 (.A(_05483_),
    .X(net269));
 sky130_fd_sc_hd__buf_12 max_cap270 (.A(_05481_),
    .X(net270));
 sky130_fd_sc_hd__buf_12 max_cap271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_12 max_cap272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_12 max_cap273 (.A(_05233_),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_16 max_cap274 (.A(_05233_),
    .X(net274));
 sky130_fd_sc_hd__buf_12 max_cap275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__buf_12 max_cap276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_12 max_cap277 (.A(_04029_),
    .X(net277));
 sky130_fd_sc_hd__buf_12 max_cap278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_12 max_cap279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_12 max_cap280 (.A(_01962_),
    .X(net280));
 sky130_fd_sc_hd__buf_8 max_cap281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_8 max_cap282 (.A(_06307_),
    .X(net282));
 sky130_fd_sc_hd__buf_8 max_cap283 (.A(_06307_),
    .X(net283));
 sky130_fd_sc_hd__buf_12 max_cap284 (.A(_06305_),
    .X(net284));
 sky130_fd_sc_hd__buf_8 max_cap285 (.A(_06011_),
    .X(net285));
 sky130_fd_sc_hd__buf_12 max_cap286 (.A(_06011_),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_8 max_cap287 (.A(_06010_),
    .X(net287));
 sky130_fd_sc_hd__buf_6 max_cap288 (.A(_05766_),
    .X(net288));
 sky130_fd_sc_hd__buf_12 max_cap289 (.A(_05766_),
    .X(net289));
 sky130_fd_sc_hd__buf_12 max_cap290 (.A(_05762_),
    .X(net290));
 sky130_fd_sc_hd__buf_12 max_cap291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_12 max_cap292 (.A(_05508_),
    .X(net292));
 sky130_fd_sc_hd__buf_12 wire293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__buf_12 wire294 (.A(_05249_),
    .X(net294));
 sky130_fd_sc_hd__buf_12 max_cap295 (.A(_05248_),
    .X(net295));
 sky130_fd_sc_hd__buf_8 max_cap296 (.A(_05231_),
    .X(net296));
 sky130_fd_sc_hd__buf_12 max_cap297 (.A(_05231_),
    .X(net297));
 sky130_fd_sc_hd__buf_12 max_cap298 (.A(_04238_),
    .X(net298));
 sky130_fd_sc_hd__buf_12 max_cap299 (.A(_04227_),
    .X(net299));
 sky130_fd_sc_hd__buf_12 max_cap300 (.A(_04019_),
    .X(net300));
 sky130_fd_sc_hd__buf_8 max_cap301 (.A(_04008_),
    .X(net301));
 sky130_fd_sc_hd__buf_8 max_cap302 (.A(_04008_),
    .X(net302));
 sky130_fd_sc_hd__buf_12 max_cap303 (.A(_01951_),
    .X(net303));
 sky130_fd_sc_hd__buf_8 max_cap304 (.A(_01940_),
    .X(net304));
 sky130_fd_sc_hd__buf_6 max_cap305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_8 max_cap306 (.A(_01940_),
    .X(net306));
 sky130_fd_sc_hd__buf_12 max_cap307 (.A(net309),
    .X(net307));
 sky130_fd_sc_hd__buf_12 max_cap308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__buf_12 max_cap309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__buf_12 max_cap310 (.A(_00055_),
    .X(net310));
 sky130_fd_sc_hd__buf_12 max_cap311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__buf_12 max_cap312 (.A(net313),
    .X(net312));
 sky130_fd_sc_hd__buf_12 max_cap313 (.A(_12692_),
    .X(net313));
 sky130_fd_sc_hd__buf_8 max_cap314 (.A(net317),
    .X(net314));
 sky130_fd_sc_hd__buf_8 max_cap315 (.A(net316),
    .X(net315));
 sky130_fd_sc_hd__buf_8 max_cap316 (.A(_05244_),
    .X(net316));
 sky130_fd_sc_hd__buf_6 max_cap317 (.A(_05244_),
    .X(net317));
 sky130_fd_sc_hd__buf_12 max_cap318 (.A(_05242_),
    .X(net318));
 sky130_fd_sc_hd__buf_12 max_cap319 (.A(_00251_),
    .X(net319));
 sky130_fd_sc_hd__buf_12 wire320 (.A(_00240_),
    .X(net320));
 sky130_fd_sc_hd__buf_6 max_cap321 (.A(net323),
    .X(net321));
 sky130_fd_sc_hd__buf_8 max_cap322 (.A(_00033_),
    .X(net322));
 sky130_fd_sc_hd__buf_12 max_cap323 (.A(_00033_),
    .X(net323));
 sky130_fd_sc_hd__buf_12 max_cap324 (.A(_00011_),
    .X(net324));
 sky130_fd_sc_hd__buf_12 max_cap325 (.A(net326),
    .X(net325));
 sky130_fd_sc_hd__buf_12 max_cap326 (.A(_12899_),
    .X(net326));
 sky130_fd_sc_hd__buf_12 max_cap327 (.A(_12681_),
    .X(net327));
 sky130_fd_sc_hd__buf_8 max_cap328 (.A(_12670_),
    .X(net328));
 sky130_fd_sc_hd__buf_8 max_cap329 (.A(_12670_),
    .X(net329));
 sky130_fd_sc_hd__buf_12 wire330 (.A(_11309_),
    .X(net330));
 sky130_fd_sc_hd__buf_12 wire331 (.A(_11298_),
    .X(net331));
 sky130_fd_sc_hd__buf_12 max_cap332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__buf_12 max_cap333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__buf_12 max_cap334 (.A(_11068_),
    .X(net334));
 sky130_fd_sc_hd__buf_12 max_cap335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__buf_12 max_cap336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_12 max_cap337 (.A(_09829_),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_16 max_cap338 (.A(_08721_),
    .X(net338));
 sky130_fd_sc_hd__buf_4 max_cap339 (.A(_04161_),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_8 max_cap340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__buf_4 max_cap341 (.A(_04161_),
    .X(net341));
 sky130_fd_sc_hd__buf_8 wire342 (.A(_02071_),
    .X(net342));
 sky130_fd_sc_hd__buf_8 max_cap343 (.A(_02071_),
    .X(net343));
 sky130_fd_sc_hd__buf_12 max_cap344 (.A(_00196_),
    .X(net344));
 sky130_fd_sc_hd__buf_12 max_cap345 (.A(_12856_),
    .X(net345));
 sky130_fd_sc_hd__buf_12 max_cap346 (.A(_11057_),
    .X(net346));
 sky130_fd_sc_hd__buf_12 max_cap347 (.A(_11046_),
    .X(net347));
 sky130_fd_sc_hd__buf_12 wire348 (.A(_10025_),
    .X(net348));
 sky130_fd_sc_hd__buf_12 max_cap349 (.A(_09807_),
    .X(net349));
 sky130_fd_sc_hd__buf_8 max_cap350 (.A(_09785_),
    .X(net350));
 sky130_fd_sc_hd__buf_8 max_cap351 (.A(_09785_),
    .X(net351));
 sky130_fd_sc_hd__buf_12 max_cap352 (.A(_08700_),
    .X(net352));
 sky130_fd_sc_hd__buf_12 max_cap353 (.A(_08678_),
    .X(net353));
 sky130_fd_sc_hd__buf_12 max_cap354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__buf_12 max_cap355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__buf_12 max_cap356 (.A(_07713_),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_16 max_cap357 (.A(_06837_),
    .X(net357));
 sky130_fd_sc_hd__buf_12 max_cap358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_12 wire359 (.A(_05720_),
    .X(net359));
 sky130_fd_sc_hd__buf_12 max_cap360 (.A(_05720_),
    .X(net360));
 sky130_fd_sc_hd__buf_12 max_cap361 (.A(_12845_),
    .X(net361));
 sky130_fd_sc_hd__buf_8 max_cap362 (.A(net364),
    .X(net362));
 sky130_fd_sc_hd__buf_8 max_cap363 (.A(_09993_),
    .X(net363));
 sky130_fd_sc_hd__buf_8 max_cap364 (.A(_09993_),
    .X(net364));
 sky130_fd_sc_hd__buf_12 max_cap365 (.A(_09971_),
    .X(net365));
 sky130_fd_sc_hd__buf_12 max_cap366 (.A(_08885_),
    .X(net366));
 sky130_fd_sc_hd__buf_12 max_cap367 (.A(_08841_),
    .X(net367));
 sky130_fd_sc_hd__buf_8 max_cap368 (.A(_07844_),
    .X(net368));
 sky130_fd_sc_hd__buf_8 max_cap369 (.A(_07844_),
    .X(net369));
 sky130_fd_sc_hd__buf_6 max_cap370 (.A(_07822_),
    .X(net370));
 sky130_fd_sc_hd__buf_12 max_cap371 (.A(_07702_),
    .X(net371));
 sky130_fd_sc_hd__buf_8 max_cap372 (.A(net373),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_8 max_cap373 (.A(_07691_),
    .X(net373));
 sky130_fd_sc_hd__buf_12 max_cap374 (.A(_07691_),
    .X(net374));
 sky130_fd_sc_hd__buf_8 max_cap375 (.A(_07011_),
    .X(net375));
 sky130_fd_sc_hd__buf_6 max_cap376 (.A(_07000_),
    .X(net376));
 sky130_fd_sc_hd__buf_8 max_cap377 (.A(_06967_),
    .X(net377));
 sky130_fd_sc_hd__buf_12 max_cap378 (.A(_06815_),
    .X(net378));
 sky130_fd_sc_hd__buf_12 max_cap379 (.A(_06793_),
    .X(net379));
 sky130_fd_sc_hd__buf_8 max_cap380 (.A(_06289_),
    .X(net380));
 sky130_fd_sc_hd__buf_8 max_cap381 (.A(_06289_),
    .X(net381));
 sky130_fd_sc_hd__buf_8 max_cap382 (.A(_06267_),
    .X(net382));
 sky130_fd_sc_hd__buf_12 max_cap383 (.A(_05698_),
    .X(net383));
 sky130_fd_sc_hd__buf_12 max_cap384 (.A(_05676_),
    .X(net384));
 sky130_fd_sc_hd__buf_8 max_cap385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_8 max_cap386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__buf_8 max_cap387 (.A(_05545_),
    .X(net387));
 sky130_fd_sc_hd__buf_12 max_cap388 (.A(_05403_),
    .X(net388));
 sky130_fd_sc_hd__buf_4 max_cap389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__buf_4 max_cap390 (.A(_07800_),
    .X(net390));
 sky130_fd_sc_hd__buf_12 max_cap391 (.A(_06310_),
    .X(net391));
 sky130_fd_sc_hd__buf_4 max_cap392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_8 max_cap393 (.A(_06245_),
    .X(net393));
 sky130_fd_sc_hd__buf_4 max_cap394 (.A(_06245_),
    .X(net394));
 sky130_fd_sc_hd__buf_6 max_cap395 (.A(_05774_),
    .X(net395));
 sky130_fd_sc_hd__buf_12 max_cap396 (.A(_05534_),
    .X(net396));
 sky130_fd_sc_hd__buf_12 max_cap397 (.A(_05469_),
    .X(net397));
 sky130_fd_sc_hd__buf_12 max_cap398 (.A(_05447_),
    .X(net398));
 sky130_fd_sc_hd__buf_8 max_cap399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__buf_8 max_cap400 (.A(_05370_),
    .X(net400));
 sky130_fd_sc_hd__buf_8 max_cap401 (.A(_05370_),
    .X(net401));
 sky130_fd_sc_hd__buf_12 max_cap402 (.A(_05348_),
    .X(net402));
 sky130_fd_sc_hd__buf_12 max_cap403 (.A(_05239_),
    .X(net403));
 sky130_fd_sc_hd__buf_12 max_cap404 (.A(_05174_),
    .X(net404));
 sky130_fd_sc_hd__buf_12 max_cap405 (.A(_05174_),
    .X(net405));
 sky130_fd_sc_hd__buf_4 max_cap406 (.A(_05818_),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_8 max_cap407 (.A(_05196_),
    .X(net407));
 sky130_fd_sc_hd__buf_12 max_cap408 (.A(_05130_),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_16 max_cap409 (.A(net57),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_16 max_cap410 (.A(net25),
    .X(net410));
endmodule
