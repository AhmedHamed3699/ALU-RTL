module CarryBypassAdder (Cin,
    Cout,
    Overflow,
    A,
    B,
    Sum);
 input Cin;
 output Cout;
 output Overflow;
 input [31:0] A;
 input [31:0] B;
 output [31:0] Sum;

 wire \BLOCKS[0].ADDERS[0].genblk1.FA.sum ;
 wire \BLOCKS[0].ADDERS[1].genblk1.FA.sum ;
 wire \BLOCKS[0].ADDERS[2].genblk1.FA.sum ;
 wire \BLOCKS[0].ADDERS[3].genblk1.FA.sum ;
 wire \BLOCKS[1].ADDERS[0].genblk1.FA.sum ;
 wire \BLOCKS[1].ADDERS[1].genblk1.FA.sum ;
 wire \BLOCKS[1].ADDERS[2].genblk1.FA.sum ;
 wire \BLOCKS[1].ADDERS[3].genblk1.FA.sum ;
 wire \BLOCKS[2].ADDERS[0].genblk1.FA.sum ;
 wire \BLOCKS[2].ADDERS[1].genblk1.FA.sum ;
 wire \BLOCKS[2].ADDERS[2].genblk1.FA.sum ;
 wire \BLOCKS[2].ADDERS[3].genblk1.FA.sum ;
 wire \BLOCKS[3].ADDERS[0].genblk1.FA.sum ;
 wire \BLOCKS[3].ADDERS[1].genblk1.FA.sum ;
 wire \BLOCKS[3].ADDERS[2].genblk1.FA.sum ;
 wire \BLOCKS[3].ADDERS[3].genblk1.FA.sum ;
 wire \BLOCKS[4].ADDERS[0].genblk1.FA.sum ;
 wire \BLOCKS[4].ADDERS[1].genblk1.FA.sum ;
 wire \BLOCKS[4].ADDERS[2].genblk1.FA.sum ;
 wire \BLOCKS[4].ADDERS[3].genblk1.FA.sum ;
 wire \BLOCKS[5].ADDERS[0].genblk1.FA.sum ;
 wire \BLOCKS[5].ADDERS[1].genblk1.FA.sum ;
 wire \BLOCKS[5].ADDERS[2].genblk1.FA.sum ;
 wire \BLOCKS[5].ADDERS[3].genblk1.FA.sum ;
 wire \BLOCKS[6].ADDERS[0].genblk1.FA.sum ;
 wire \BLOCKS[6].ADDERS[1].genblk1.FA.sum ;
 wire \BLOCKS[6].ADDERS[2].genblk1.FA.sum ;
 wire \BLOCKS[6].ADDERS[3].genblk1.FA.sum ;
 wire \BLOCKS[7].ADDERS[0].genblk1.FA.sum ;
 wire \BLOCKS[7].ADDERS[1].genblk1.FA.sum ;
 wire \BLOCKS[7].ADDERS[2].genblk1.FA.sum ;
 wire \BLOCKS[7].ADDERS[3].genblk1.FA.sum ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__inv_2 _231_ (.A(net54),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _232_ (.A(net22),
    .Y(_001_));
 sky130_fd_sc_hd__and2b_1 _233_ (.A_N(net57),
    .B(net25),
    .X(_002_));
 sky130_fd_sc_hd__and2b_1 _234_ (.A_N(net25),
    .B(net57),
    .X(_003_));
 sky130_fd_sc_hd__nor2_1 _235_ (.A(_002_),
    .B(_003_),
    .Y(_004_));
 sky130_fd_sc_hd__nand2_1 _236_ (.A(net56),
    .B(net24),
    .Y(_005_));
 sky130_fd_sc_hd__and2b_1 _237_ (.A_N(net56),
    .B(net24),
    .X(_006_));
 sky130_fd_sc_hd__and2b_1 _238_ (.A_N(net24),
    .B(net56),
    .X(_007_));
 sky130_fd_sc_hd__or2_1 _239_ (.A(_006_),
    .B(_007_),
    .X(_008_));
 sky130_fd_sc_hd__nor2_1 _240_ (.A(_000_),
    .B(_001_),
    .Y(_009_));
 sky130_fd_sc_hd__nor2_1 _241_ (.A(net54),
    .B(_001_),
    .Y(_010_));
 sky130_fd_sc_hd__nor2_1 _242_ (.A(net22),
    .B(_000_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_1 _243_ (.A(_010_),
    .B(_011_),
    .Y(_012_));
 sky130_fd_sc_hd__and2_1 _244_ (.A(net53),
    .B(net21),
    .X(_013_));
 sky130_fd_sc_hd__nand2_1 _245_ (.A(net53),
    .B(net21),
    .Y(_014_));
 sky130_fd_sc_hd__and2b_1 _246_ (.A_N(net52),
    .B(net20),
    .X(_015_));
 sky130_fd_sc_hd__and2b_1 _247_ (.A_N(net20),
    .B(net52),
    .X(_016_));
 sky130_fd_sc_hd__nor2_1 _248_ (.A(_015_),
    .B(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__and2_1 _249_ (.A(net51),
    .B(net19),
    .X(_018_));
 sky130_fd_sc_hd__nand2_1 _250_ (.A(net51),
    .B(net19),
    .Y(_019_));
 sky130_fd_sc_hd__and2b_1 _251_ (.A_N(net51),
    .B(net19),
    .X(_020_));
 sky130_fd_sc_hd__and2b_1 _252_ (.A_N(net19),
    .B(net51),
    .X(_021_));
 sky130_fd_sc_hd__nor2_1 _253_ (.A(_020_),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__and2_1 _254_ (.A(net50),
    .B(net18),
    .X(_023_));
 sky130_fd_sc_hd__nand2_1 _255_ (.A(net50),
    .B(net18),
    .Y(_024_));
 sky130_fd_sc_hd__and2b_1 _256_ (.A_N(net50),
    .B(net18),
    .X(_025_));
 sky130_fd_sc_hd__and2b_1 _257_ (.A_N(net18),
    .B(net50),
    .X(_026_));
 sky130_fd_sc_hd__nor2_1 _258_ (.A(_025_),
    .B(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__and2_1 _259_ (.A(net49),
    .B(net17),
    .X(_028_));
 sky130_fd_sc_hd__nand2_1 _260_ (.A(net49),
    .B(net17),
    .Y(_029_));
 sky130_fd_sc_hd__and2b_1 _261_ (.A_N(net48),
    .B(net16),
    .X(_030_));
 sky130_fd_sc_hd__and2b_1 _262_ (.A_N(net16),
    .B(net48),
    .X(_031_));
 sky130_fd_sc_hd__and2_1 _263_ (.A(net47),
    .B(net15),
    .X(_032_));
 sky130_fd_sc_hd__nand2_1 _264_ (.A(net47),
    .B(net15),
    .Y(_033_));
 sky130_fd_sc_hd__and2b_1 _265_ (.A_N(net47),
    .B(net15),
    .X(_034_));
 sky130_fd_sc_hd__and2b_1 _266_ (.A_N(net15),
    .B(net47),
    .X(_035_));
 sky130_fd_sc_hd__nor2_1 _267_ (.A(_034_),
    .B(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__and2_1 _268_ (.A(net46),
    .B(net14),
    .X(_037_));
 sky130_fd_sc_hd__nand2_1 _269_ (.A(net46),
    .B(net14),
    .Y(_038_));
 sky130_fd_sc_hd__and2b_1 _270_ (.A_N(net46),
    .B(net14),
    .X(_039_));
 sky130_fd_sc_hd__and2b_1 _271_ (.A_N(net14),
    .B(net46),
    .X(_040_));
 sky130_fd_sc_hd__and2_1 _272_ (.A(net45),
    .B(net13),
    .X(_041_));
 sky130_fd_sc_hd__nand2_1 _273_ (.A(net45),
    .B(net13),
    .Y(_042_));
 sky130_fd_sc_hd__and2b_1 _274_ (.A_N(net43),
    .B(net11),
    .X(_043_));
 sky130_fd_sc_hd__and2b_1 _275_ (.A_N(net11),
    .B(net43),
    .X(_044_));
 sky130_fd_sc_hd__and2_1 _276_ (.A(net42),
    .B(net10),
    .X(_045_));
 sky130_fd_sc_hd__nand2_1 _277_ (.A(net42),
    .B(net10),
    .Y(_046_));
 sky130_fd_sc_hd__and2b_1 _278_ (.A_N(net42),
    .B(net10),
    .X(_047_));
 sky130_fd_sc_hd__and2b_1 _279_ (.A_N(net10),
    .B(net42),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _280_ (.A(net41),
    .B(net9),
    .X(_049_));
 sky130_fd_sc_hd__nand2_1 _281_ (.A(net41),
    .B(net9),
    .Y(_050_));
 sky130_fd_sc_hd__or2_1 _282_ (.A(net41),
    .B(net9),
    .X(_051_));
 sky130_fd_sc_hd__and2b_1 _283_ (.A_N(net41),
    .B(net9),
    .X(_052_));
 sky130_fd_sc_hd__and2b_1 _284_ (.A_N(net9),
    .B(net41),
    .X(_053_));
 sky130_fd_sc_hd__and2_1 _285_ (.A(net40),
    .B(net8),
    .X(_054_));
 sky130_fd_sc_hd__nand2_1 _286_ (.A(net40),
    .B(net8),
    .Y(_055_));
 sky130_fd_sc_hd__and2b_1 _287_ (.A_N(net39),
    .B(net7),
    .X(_056_));
 sky130_fd_sc_hd__and2b_1 _288_ (.A_N(net7),
    .B(net39),
    .X(_057_));
 sky130_fd_sc_hd__nor2_1 _289_ (.A(_056_),
    .B(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__and2_1 _290_ (.A(net38),
    .B(net6),
    .X(_059_));
 sky130_fd_sc_hd__nand2_1 _291_ (.A(net38),
    .B(net6),
    .Y(_060_));
 sky130_fd_sc_hd__and2b_1 _292_ (.A_N(net38),
    .B(net6),
    .X(_061_));
 sky130_fd_sc_hd__and2b_1 _293_ (.A_N(net6),
    .B(net38),
    .X(_062_));
 sky130_fd_sc_hd__nor2_1 _294_ (.A(_061_),
    .B(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__and2_1 _295_ (.A(net37),
    .B(net5),
    .X(_064_));
 sky130_fd_sc_hd__nand2_1 _296_ (.A(net37),
    .B(net5),
    .Y(_065_));
 sky130_fd_sc_hd__and2b_1 _297_ (.A_N(net37),
    .B(net5),
    .X(_066_));
 sky130_fd_sc_hd__and2b_1 _298_ (.A_N(net5),
    .B(net37),
    .X(_067_));
 sky130_fd_sc_hd__nor2_1 _299_ (.A(_066_),
    .B(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__and2_1 _300_ (.A(net36),
    .B(net4),
    .X(_069_));
 sky130_fd_sc_hd__nand2_1 _301_ (.A(net36),
    .B(net4),
    .Y(_070_));
 sky130_fd_sc_hd__and2_1 _302_ (.A(net34),
    .B(net2),
    .X(_071_));
 sky130_fd_sc_hd__nand2_1 _303_ (.A(net34),
    .B(net2),
    .Y(_072_));
 sky130_fd_sc_hd__and2_1 _304_ (.A(net64),
    .B(net32),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _305_ (.A(net63),
    .B(net31),
    .X(_074_));
 sky130_fd_sc_hd__and2_1 _306_ (.A(net62),
    .B(net30),
    .X(_075_));
 sky130_fd_sc_hd__and2_1 _307_ (.A(net61),
    .B(net29),
    .X(_076_));
 sky130_fd_sc_hd__nor2_1 _308_ (.A(net61),
    .B(net29),
    .Y(_077_));
 sky130_fd_sc_hd__nor2_1 _309_ (.A(_076_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__and2_1 _310_ (.A(net60),
    .B(net28),
    .X(_079_));
 sky130_fd_sc_hd__and2_1 _311_ (.A(net59),
    .B(net27),
    .X(_080_));
 sky130_fd_sc_hd__nor2_1 _312_ (.A(net59),
    .B(net27),
    .Y(_081_));
 sky130_fd_sc_hd__nor2_1 _313_ (.A(_080_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__and2_1 _314_ (.A(net58),
    .B(net26),
    .X(_083_));
 sky130_fd_sc_hd__and2_1 _315_ (.A(net55),
    .B(net23),
    .X(_084_));
 sky130_fd_sc_hd__nand2_1 _316_ (.A(net55),
    .B(net23),
    .Y(_085_));
 sky130_fd_sc_hd__or2_1 _317_ (.A(net55),
    .B(net23),
    .X(_086_));
 sky130_fd_sc_hd__or2_1 _318_ (.A(net44),
    .B(net12),
    .X(_087_));
 sky130_fd_sc_hd__nand2_1 _319_ (.A(net44),
    .B(net12),
    .Y(_088_));
 sky130_fd_sc_hd__or2_1 _320_ (.A(net33),
    .B(net1),
    .X(_089_));
 sky130_fd_sc_hd__nand2_1 _321_ (.A(net33),
    .B(net1),
    .Y(_090_));
 sky130_fd_sc_hd__o21ai_1 _322_ (.A1(net33),
    .A2(net1),
    .B1(net65),
    .Y(_091_));
 sky130_fd_sc_hd__and2_1 _323_ (.A(_090_),
    .B(_091_),
    .X(_092_));
 sky130_fd_sc_hd__nand3_1 _324_ (.A(_088_),
    .B(_090_),
    .C(_091_),
    .Y(_093_));
 sky130_fd_sc_hd__o21a_1 _325_ (.A1(net44),
    .A2(net12),
    .B1(_093_),
    .X(_094_));
 sky130_fd_sc_hd__and3_1 _326_ (.A(_094_),
    .B(_086_),
    .C(_085_),
    .X(_095_));
 sky130_fd_sc_hd__a31oi_2 _327_ (.A1(_086_),
    .A2(_087_),
    .A3(_093_),
    .B1(_084_),
    .Y(_096_));
 sky130_fd_sc_hd__nor2_1 _328_ (.A(net58),
    .B(net26),
    .Y(_097_));
 sky130_fd_sc_hd__or2_1 _329_ (.A(_083_),
    .B(_097_),
    .X(_098_));
 sky130_fd_sc_hd__o21bai_1 _330_ (.A1(_098_),
    .A2(_096_),
    .B1_N(_083_),
    .Y(_099_));
 sky130_fd_sc_hd__a21oi_1 _331_ (.A1(_099_),
    .A2(_082_),
    .B1(_080_),
    .Y(_100_));
 sky130_fd_sc_hd__nor2_1 _332_ (.A(net60),
    .B(net28),
    .Y(_101_));
 sky130_fd_sc_hd__or2_1 _333_ (.A(_079_),
    .B(_101_),
    .X(_102_));
 sky130_fd_sc_hd__o21bai_1 _334_ (.A1(_102_),
    .A2(_100_),
    .B1_N(_079_),
    .Y(_103_));
 sky130_fd_sc_hd__a21oi_1 _335_ (.A1(_103_),
    .A2(_078_),
    .B1(_076_),
    .Y(_104_));
 sky130_fd_sc_hd__nor2_1 _336_ (.A(net62),
    .B(net30),
    .Y(_105_));
 sky130_fd_sc_hd__or2_1 _337_ (.A(_075_),
    .B(_105_),
    .X(_106_));
 sky130_fd_sc_hd__o21bai_1 _338_ (.A1(_106_),
    .A2(_104_),
    .B1_N(_075_),
    .Y(_107_));
 sky130_fd_sc_hd__or2_1 _339_ (.A(net63),
    .B(net31),
    .X(_108_));
 sky130_fd_sc_hd__nand2b_1 _340_ (.A_N(_074_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__a21oi_1 _341_ (.A1(_107_),
    .A2(_108_),
    .B1(_074_),
    .Y(_110_));
 sky130_fd_sc_hd__nor2_1 _342_ (.A(net64),
    .B(net32),
    .Y(_111_));
 sky130_fd_sc_hd__or2_1 _343_ (.A(_073_),
    .B(_111_),
    .X(_112_));
 sky130_fd_sc_hd__o21bai_2 _344_ (.A1(_112_),
    .A2(_110_),
    .B1_N(_073_),
    .Y(_113_));
 sky130_fd_sc_hd__or2_1 _345_ (.A(net34),
    .B(net2),
    .X(_114_));
 sky130_fd_sc_hd__nand2_1 _346_ (.A(_072_),
    .B(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _347_ (.A(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__nand2_1 _348_ (.A(_113_),
    .B(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__a21oi_1 _349_ (.A1(_113_),
    .A2(_116_),
    .B1(_071_),
    .Y(_118_));
 sky130_fd_sc_hd__and2b_1 _350_ (.A_N(net35),
    .B(net3),
    .X(_119_));
 sky130_fd_sc_hd__and2b_1 _351_ (.A_N(net3),
    .B(net35),
    .X(_120_));
 sky130_fd_sc_hd__nor2_1 _352_ (.A(_119_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__o2bb2ai_1 _353_ (.A1_N(_072_),
    .A2_N(_117_),
    .B1(_119_),
    .B2(_120_),
    .Y(_122_));
 sky130_fd_sc_hd__or4_1 _354_ (.A(_109_),
    .B(_112_),
    .C(_115_),
    .D(_121_),
    .X(_123_));
 sky130_fd_sc_hd__a21bo_1 _355_ (.A1(net35),
    .A2(net3),
    .B1_N(_123_),
    .X(_124_));
 sky130_fd_sc_hd__inv_2 _356_ (.A(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__o21bai_2 _357_ (.A1(_121_),
    .A2(_118_),
    .B1_N(_124_),
    .Y(_126_));
 sky130_fd_sc_hd__or2_1 _358_ (.A(net36),
    .B(net4),
    .X(_127_));
 sky130_fd_sc_hd__or2_1 _359_ (.A(_107_),
    .B(_123_),
    .X(_128_));
 sky130_fd_sc_hd__nand2_1 _360_ (.A(_070_),
    .B(_127_),
    .Y(_129_));
 sky130_fd_sc_hd__and3_1 _361_ (.A(_070_),
    .B(_127_),
    .C(_128_),
    .X(_130_));
 sky130_fd_sc_hd__a21boi_1 _362_ (.A1(_122_),
    .A2(_125_),
    .B1_N(_130_),
    .Y(_131_));
 sky130_fd_sc_hd__nand2_1 _363_ (.A(_126_),
    .B(_130_),
    .Y(_132_));
 sky130_fd_sc_hd__a2bb2oi_1 _364_ (.A1_N(_066_),
    .A2_N(_067_),
    .B1(_070_),
    .B2(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__o22ai_1 _365_ (.A1(_066_),
    .A2(_067_),
    .B1(_069_),
    .B2(_131_),
    .Y(_134_));
 sky130_fd_sc_hd__a2bb2oi_1 _366_ (.A1_N(_061_),
    .A2_N(_062_),
    .B1(_065_),
    .B2(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__o22ai_1 _367_ (.A1(_061_),
    .A2(_062_),
    .B1(_064_),
    .B2(_133_),
    .Y(_136_));
 sky130_fd_sc_hd__a2bb2oi_1 _368_ (.A1_N(_056_),
    .A2_N(_057_),
    .B1(_060_),
    .B2(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__o22ai_1 _369_ (.A1(_056_),
    .A2(_057_),
    .B1(_059_),
    .B2(_135_),
    .Y(_138_));
 sky130_fd_sc_hd__or4_1 _370_ (.A(_058_),
    .B(_063_),
    .C(_068_),
    .D(_129_),
    .X(_139_));
 sky130_fd_sc_hd__a21boi_2 _371_ (.A1(net39),
    .A2(net7),
    .B1_N(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__inv_2 _372_ (.A(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__or2_1 _373_ (.A(net40),
    .B(net8),
    .X(_142_));
 sky130_fd_sc_hd__a21oi_1 _374_ (.A1(_126_),
    .A2(_128_),
    .B1(_139_),
    .Y(_143_));
 sky130_fd_sc_hd__nand2_1 _375_ (.A(_055_),
    .B(_142_),
    .Y(_144_));
 sky130_fd_sc_hd__or2_1 _376_ (.A(_144_),
    .B(_143_),
    .X(_145_));
 sky130_fd_sc_hd__a21oi_1 _377_ (.A1(_138_),
    .A2(_140_),
    .B1(_143_),
    .Y(_146_));
 sky130_fd_sc_hd__a21oi_1 _378_ (.A1(_138_),
    .A2(_140_),
    .B1(_145_),
    .Y(_147_));
 sky130_fd_sc_hd__o21bai_1 _379_ (.A1(_141_),
    .A2(_137_),
    .B1_N(_145_),
    .Y(_148_));
 sky130_fd_sc_hd__a2bb2oi_1 _380_ (.A1_N(_052_),
    .A2_N(_053_),
    .B1(_055_),
    .B2(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__o22ai_1 _381_ (.A1(_052_),
    .A2(_053_),
    .B1(_054_),
    .B2(_147_),
    .Y(_150_));
 sky130_fd_sc_hd__a2bb2oi_1 _382_ (.A1_N(_047_),
    .A2_N(_048_),
    .B1(_050_),
    .B2(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__o22ai_1 _383_ (.A1(_047_),
    .A2(_048_),
    .B1(_049_),
    .B2(_149_),
    .Y(_152_));
 sky130_fd_sc_hd__a2bb2oi_1 _384_ (.A1_N(_043_),
    .A2_N(_044_),
    .B1(_046_),
    .B2(_152_),
    .Y(_153_));
 sky130_fd_sc_hd__o22ai_1 _385_ (.A1(_043_),
    .A2(_044_),
    .B1(_045_),
    .B2(_151_),
    .Y(_154_));
 sky130_fd_sc_hd__o22a_1 _386_ (.A1(_043_),
    .A2(_044_),
    .B1(_047_),
    .B2(_048_),
    .X(_155_));
 sky130_fd_sc_hd__or4bb_1 _387_ (.A(_049_),
    .B(_144_),
    .C_N(_155_),
    .D_N(_051_),
    .X(_156_));
 sky130_fd_sc_hd__a21boi_1 _388_ (.A1(net43),
    .A2(net11),
    .B1_N(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__a21bo_1 _389_ (.A1(net43),
    .A2(net11),
    .B1_N(_156_),
    .X(_158_));
 sky130_fd_sc_hd__nor2_1 _390_ (.A(net45),
    .B(net13),
    .Y(_159_));
 sky130_fd_sc_hd__nor2_1 _391_ (.A(_041_),
    .B(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__o21ai_1 _392_ (.A1(_156_),
    .A2(_146_),
    .B1(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__o22a_1 _393_ (.A1(_146_),
    .A2(_156_),
    .B1(_158_),
    .B2(_153_),
    .X(_162_));
 sky130_fd_sc_hd__a21oi_1 _394_ (.A1(_154_),
    .A2(_157_),
    .B1(_161_),
    .Y(_163_));
 sky130_fd_sc_hd__o21bai_1 _395_ (.A1(_158_),
    .A2(_153_),
    .B1_N(_161_),
    .Y(_164_));
 sky130_fd_sc_hd__a2bb2oi_1 _396_ (.A1_N(_039_),
    .A2_N(_040_),
    .B1(_042_),
    .B2(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__o22ai_1 _397_ (.A1(_039_),
    .A2(_040_),
    .B1(_041_),
    .B2(_163_),
    .Y(_166_));
 sky130_fd_sc_hd__a2bb2oi_1 _398_ (.A1_N(_034_),
    .A2_N(_035_),
    .B1(_038_),
    .B2(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__o22ai_1 _399_ (.A1(_034_),
    .A2(_035_),
    .B1(_037_),
    .B2(_165_),
    .Y(_168_));
 sky130_fd_sc_hd__a2bb2oi_1 _400_ (.A1_N(_030_),
    .A2_N(_031_),
    .B1(_033_),
    .B2(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__o22ai_1 _401_ (.A1(_030_),
    .A2(_031_),
    .B1(_032_),
    .B2(_167_),
    .Y(_170_));
 sky130_fd_sc_hd__o22a_1 _402_ (.A1(_030_),
    .A2(_031_),
    .B1(_034_),
    .B2(_035_),
    .X(_171_));
 sky130_fd_sc_hd__o211ai_2 _403_ (.A1(_039_),
    .A2(_040_),
    .B1(_160_),
    .C1(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__a21boi_1 _404_ (.A1(net48),
    .A2(net16),
    .B1_N(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__inv_2 _405_ (.A(_173_),
    .Y(_174_));
 sky130_fd_sc_hd__or2_1 _406_ (.A(net49),
    .B(net17),
    .X(_175_));
 sky130_fd_sc_hd__nand2_1 _407_ (.A(_029_),
    .B(_175_),
    .Y(_176_));
 sky130_fd_sc_hd__o211ai_1 _408_ (.A1(_172_),
    .A2(_162_),
    .B1(_029_),
    .C1(_175_),
    .Y(_177_));
 sky130_fd_sc_hd__o22a_1 _409_ (.A1(_162_),
    .A2(_172_),
    .B1(_174_),
    .B2(_169_),
    .X(_178_));
 sky130_fd_sc_hd__a21oi_1 _410_ (.A1(_170_),
    .A2(_173_),
    .B1(_177_),
    .Y(_179_));
 sky130_fd_sc_hd__o21bai_1 _411_ (.A1(_174_),
    .A2(_169_),
    .B1_N(_177_),
    .Y(_180_));
 sky130_fd_sc_hd__a2bb2oi_1 _412_ (.A1_N(_025_),
    .A2_N(_026_),
    .B1(_029_),
    .B2(_180_),
    .Y(_181_));
 sky130_fd_sc_hd__o22ai_1 _413_ (.A1(_025_),
    .A2(_026_),
    .B1(_028_),
    .B2(_179_),
    .Y(_182_));
 sky130_fd_sc_hd__a21oi_1 _414_ (.A1(_024_),
    .A2(_182_),
    .B1(_022_),
    .Y(_183_));
 sky130_fd_sc_hd__o22ai_1 _415_ (.A1(_020_),
    .A2(_021_),
    .B1(_023_),
    .B2(_181_),
    .Y(_184_));
 sky130_fd_sc_hd__a2bb2oi_1 _416_ (.A1_N(_015_),
    .A2_N(_016_),
    .B1(_019_),
    .B2(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__o22ai_1 _417_ (.A1(_015_),
    .A2(_016_),
    .B1(_018_),
    .B2(_183_),
    .Y(_186_));
 sky130_fd_sc_hd__or4_1 _418_ (.A(_017_),
    .B(_022_),
    .C(_027_),
    .D(_176_),
    .X(_187_));
 sky130_fd_sc_hd__a21boi_1 _419_ (.A1(net52),
    .A2(net20),
    .B1_N(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__a21bo_1 _420_ (.A1(net52),
    .A2(net20),
    .B1_N(_187_),
    .X(_189_));
 sky130_fd_sc_hd__or2_1 _421_ (.A(net53),
    .B(net21),
    .X(_190_));
 sky130_fd_sc_hd__o211ai_1 _422_ (.A1(_187_),
    .A2(_178_),
    .B1(_014_),
    .C1(_190_),
    .Y(_191_));
 sky130_fd_sc_hd__a21oi_1 _423_ (.A1(_186_),
    .A2(_188_),
    .B1(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__o21bai_1 _424_ (.A1(_189_),
    .A2(_185_),
    .B1_N(_191_),
    .Y(_193_));
 sky130_fd_sc_hd__a21o_1 _425_ (.A1(net53),
    .A2(net21),
    .B1(_192_),
    .X(_194_));
 sky130_fd_sc_hd__a2bb2oi_1 _426_ (.A1_N(_010_),
    .A2_N(_011_),
    .B1(_014_),
    .B2(_193_),
    .Y(_195_));
 sky130_fd_sc_hd__o22ai_1 _427_ (.A1(_010_),
    .A2(_011_),
    .B1(_013_),
    .B2(_192_),
    .Y(_196_));
 sky130_fd_sc_hd__o21ai_1 _428_ (.A1(_000_),
    .A2(_001_),
    .B1(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__o22ai_1 _429_ (.A1(_006_),
    .A2(_007_),
    .B1(_009_),
    .B2(_195_),
    .Y(_198_));
 sky130_fd_sc_hd__a21boi_1 _430_ (.A1(_197_),
    .A2(_008_),
    .B1_N(_005_),
    .Y(_199_));
 sky130_fd_sc_hd__a2bb2oi_1 _431_ (.A1_N(_002_),
    .A2_N(_003_),
    .B1(_005_),
    .B2(_198_),
    .Y(_200_));
 sky130_fd_sc_hd__o211a_1 _432_ (.A1(_010_),
    .A2(_011_),
    .B1(_014_),
    .C1(_190_),
    .X(_201_));
 sky130_fd_sc_hd__nand3b_1 _433_ (.A_N(_004_),
    .B(_008_),
    .C(_201_),
    .Y(_202_));
 sky130_fd_sc_hd__a21bo_1 _434_ (.A1(net57),
    .A2(net25),
    .B1_N(_202_),
    .X(_203_));
 sky130_fd_sc_hd__a2bb2o_1 _435_ (.A1_N(_178_),
    .A2_N(_187_),
    .B1(_188_),
    .B2(_186_),
    .X(_204_));
 sky130_fd_sc_hd__inv_2 _436_ (.A(_204_),
    .Y(_205_));
 sky130_fd_sc_hd__o22a_1 _437_ (.A1(_202_),
    .A2(_205_),
    .B1(_203_),
    .B2(_200_),
    .X(net66));
 sky130_fd_sc_hd__o22a_1 _438_ (.A1(net57),
    .A2(net25),
    .B1(_202_),
    .B2(_205_),
    .X(_206_));
 sky130_fd_sc_hd__o221ai_1 _439_ (.A1(_202_),
    .A2(_205_),
    .B1(_203_),
    .B2(_200_),
    .C1(_199_),
    .Y(_207_));
 sky130_fd_sc_hd__o21ai_1 _440_ (.A1(_199_),
    .A2(_206_),
    .B1(_207_),
    .Y(net67));
 sky130_fd_sc_hd__and3_1 _441_ (.A(net65),
    .B(net33),
    .C(net1),
    .X(_208_));
 sky130_fd_sc_hd__o22a_1 _442_ (.A1(net65),
    .A2(_089_),
    .B1(_208_),
    .B2(_092_),
    .X(\BLOCKS[0].ADDERS[0].genblk1.FA.sum ));
 sky130_fd_sc_hd__a21oi_1 _443_ (.A1(_087_),
    .A2(_088_),
    .B1(_092_),
    .Y(_209_));
 sky130_fd_sc_hd__a41o_1 _444_ (.A1(_087_),
    .A2(_088_),
    .A3(_090_),
    .A4(_091_),
    .B1(_209_),
    .X(\BLOCKS[0].ADDERS[1].genblk1.FA.sum ));
 sky130_fd_sc_hd__a21oi_1 _445_ (.A1(_085_),
    .A2(_086_),
    .B1(_094_),
    .Y(_210_));
 sky130_fd_sc_hd__nor2_1 _446_ (.A(_095_),
    .B(_210_),
    .Y(\BLOCKS[0].ADDERS[2].genblk1.FA.sum ));
 sky130_fd_sc_hd__xor2_1 _447_ (.A(_096_),
    .B(_098_),
    .X(\BLOCKS[0].ADDERS[3].genblk1.FA.sum ));
 sky130_fd_sc_hd__xor2_1 _448_ (.A(_082_),
    .B(_099_),
    .X(\BLOCKS[1].ADDERS[0].genblk1.FA.sum ));
 sky130_fd_sc_hd__xor2_1 _449_ (.A(_100_),
    .B(_102_),
    .X(\BLOCKS[1].ADDERS[1].genblk1.FA.sum ));
 sky130_fd_sc_hd__xor2_1 _450_ (.A(_078_),
    .B(_103_),
    .X(\BLOCKS[1].ADDERS[2].genblk1.FA.sum ));
 sky130_fd_sc_hd__xor2_1 _451_ (.A(_104_),
    .B(_106_),
    .X(\BLOCKS[1].ADDERS[3].genblk1.FA.sum ));
 sky130_fd_sc_hd__xnor2_1 _452_ (.A(_107_),
    .B(_109_),
    .Y(\BLOCKS[2].ADDERS[0].genblk1.FA.sum ));
 sky130_fd_sc_hd__xor2_1 _453_ (.A(_110_),
    .B(_112_),
    .X(\BLOCKS[2].ADDERS[1].genblk1.FA.sum ));
 sky130_fd_sc_hd__xnor2_1 _454_ (.A(_113_),
    .B(_115_),
    .Y(\BLOCKS[2].ADDERS[2].genblk1.FA.sum ));
 sky130_fd_sc_hd__a2111o_1 _455_ (.A1(_113_),
    .A2(_116_),
    .B1(_119_),
    .C1(_120_),
    .D1(_071_),
    .X(_211_));
 sky130_fd_sc_hd__and2_1 _456_ (.A(_122_),
    .B(_211_),
    .X(\BLOCKS[2].ADDERS[3].genblk1.FA.sum ));
 sky130_fd_sc_hd__a22oi_1 _457_ (.A1(_070_),
    .A2(_127_),
    .B1(_128_),
    .B2(_126_),
    .Y(_212_));
 sky130_fd_sc_hd__a21oi_1 _458_ (.A1(_126_),
    .A2(_130_),
    .B1(_212_),
    .Y(\BLOCKS[3].ADDERS[0].genblk1.FA.sum ));
 sky130_fd_sc_hd__or4_1 _459_ (.A(_066_),
    .B(_067_),
    .C(_069_),
    .D(_131_),
    .X(_213_));
 sky130_fd_sc_hd__and2_1 _460_ (.A(_134_),
    .B(_213_),
    .X(\BLOCKS[3].ADDERS[1].genblk1.FA.sum ));
 sky130_fd_sc_hd__and3_1 _461_ (.A(_063_),
    .B(_065_),
    .C(_134_),
    .X(_214_));
 sky130_fd_sc_hd__nor2_1 _462_ (.A(_135_),
    .B(_214_),
    .Y(\BLOCKS[3].ADDERS[2].genblk1.FA.sum ));
 sky130_fd_sc_hd__and3_1 _463_ (.A(_058_),
    .B(_060_),
    .C(_136_),
    .X(_215_));
 sky130_fd_sc_hd__nor2_1 _464_ (.A(_137_),
    .B(_215_),
    .Y(\BLOCKS[3].ADDERS[3].genblk1.FA.sum ));
 sky130_fd_sc_hd__xnor2_1 _465_ (.A(_144_),
    .B(_146_),
    .Y(\BLOCKS[4].ADDERS[0].genblk1.FA.sum ));
 sky130_fd_sc_hd__o211a_1 _466_ (.A1(_052_),
    .A2(_053_),
    .B1(_055_),
    .C1(_148_),
    .X(_216_));
 sky130_fd_sc_hd__o2bb2a_1 _467_ (.A1_N(_050_),
    .A2_N(_051_),
    .B1(_054_),
    .B2(_147_),
    .X(_217_));
 sky130_fd_sc_hd__or2_1 _468_ (.A(_216_),
    .B(_217_),
    .X(\BLOCKS[4].ADDERS[1].genblk1.FA.sum ));
 sky130_fd_sc_hd__or4_1 _469_ (.A(_047_),
    .B(_048_),
    .C(_049_),
    .D(_149_),
    .X(_218_));
 sky130_fd_sc_hd__and2_1 _470_ (.A(_152_),
    .B(_218_),
    .X(\BLOCKS[4].ADDERS[2].genblk1.FA.sum ));
 sky130_fd_sc_hd__or4_1 _471_ (.A(_043_),
    .B(_044_),
    .C(_045_),
    .D(_151_),
    .X(_219_));
 sky130_fd_sc_hd__and2_1 _472_ (.A(_154_),
    .B(_219_),
    .X(\BLOCKS[4].ADDERS[3].genblk1.FA.sum ));
 sky130_fd_sc_hd__nor2_1 _473_ (.A(_160_),
    .B(_162_),
    .Y(_220_));
 sky130_fd_sc_hd__nor2_1 _474_ (.A(_163_),
    .B(_220_),
    .Y(\BLOCKS[5].ADDERS[0].genblk1.FA.sum ));
 sky130_fd_sc_hd__or4_1 _475_ (.A(_039_),
    .B(_040_),
    .C(_041_),
    .D(_163_),
    .X(_221_));
 sky130_fd_sc_hd__and2_1 _476_ (.A(_166_),
    .B(_221_),
    .X(\BLOCKS[5].ADDERS[1].genblk1.FA.sum ));
 sky130_fd_sc_hd__and3_1 _477_ (.A(_036_),
    .B(_038_),
    .C(_166_),
    .X(_222_));
 sky130_fd_sc_hd__nor2_1 _478_ (.A(_167_),
    .B(_222_),
    .Y(\BLOCKS[5].ADDERS[2].genblk1.FA.sum ));
 sky130_fd_sc_hd__or4_1 _479_ (.A(_030_),
    .B(_031_),
    .C(_032_),
    .D(_167_),
    .X(_223_));
 sky130_fd_sc_hd__and2_1 _480_ (.A(_170_),
    .B(_223_),
    .X(\BLOCKS[5].ADDERS[3].genblk1.FA.sum ));
 sky130_fd_sc_hd__a21oi_1 _481_ (.A1(_029_),
    .A2(_175_),
    .B1(_178_),
    .Y(_224_));
 sky130_fd_sc_hd__nor2_1 _482_ (.A(_179_),
    .B(_224_),
    .Y(\BLOCKS[6].ADDERS[0].genblk1.FA.sum ));
 sky130_fd_sc_hd__or4_1 _483_ (.A(_025_),
    .B(_026_),
    .C(_028_),
    .D(_179_),
    .X(_225_));
 sky130_fd_sc_hd__and2_1 _484_ (.A(_182_),
    .B(_225_),
    .X(\BLOCKS[6].ADDERS[1].genblk1.FA.sum ));
 sky130_fd_sc_hd__and3_1 _485_ (.A(_022_),
    .B(_024_),
    .C(_182_),
    .X(_226_));
 sky130_fd_sc_hd__nor2_1 _486_ (.A(_183_),
    .B(_226_),
    .Y(\BLOCKS[6].ADDERS[2].genblk1.FA.sum ));
 sky130_fd_sc_hd__or4_1 _487_ (.A(_015_),
    .B(_016_),
    .C(_018_),
    .D(_183_),
    .X(_227_));
 sky130_fd_sc_hd__and2_1 _488_ (.A(_186_),
    .B(_227_),
    .X(\BLOCKS[6].ADDERS[3].genblk1.FA.sum ));
 sky130_fd_sc_hd__a21o_1 _489_ (.A1(_014_),
    .A2(_190_),
    .B1(_205_),
    .X(_228_));
 sky130_fd_sc_hd__and2_1 _490_ (.A(_193_),
    .B(_228_),
    .X(\BLOCKS[7].ADDERS[0].genblk1.FA.sum ));
 sky130_fd_sc_hd__xnor2_1 _491_ (.A(_012_),
    .B(_194_),
    .Y(\BLOCKS[7].ADDERS[1].genblk1.FA.sum ));
 sky130_fd_sc_hd__or4_1 _492_ (.A(_006_),
    .B(_007_),
    .C(_009_),
    .D(_195_),
    .X(_229_));
 sky130_fd_sc_hd__and2_1 _493_ (.A(_198_),
    .B(_229_),
    .X(\BLOCKS[7].ADDERS[2].genblk1.FA.sum ));
 sky130_fd_sc_hd__nand2_1 _494_ (.A(_199_),
    .B(_004_),
    .Y(_230_));
 sky130_fd_sc_hd__and2b_1 _495_ (.A_N(_200_),
    .B(_230_),
    .X(\BLOCKS[7].ADDERS[3].genblk1.FA.sum ));
 sky130_fd_sc_hd__clkbuf_1 _496_ (.A(\BLOCKS[0].ADDERS[0].genblk1.FA.sum ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _497_ (.A(\BLOCKS[0].ADDERS[1].genblk1.FA.sum ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _498_ (.A(\BLOCKS[0].ADDERS[2].genblk1.FA.sum ),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _499_ (.A(\BLOCKS[0].ADDERS[3].genblk1.FA.sum ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _500_ (.A(\BLOCKS[1].ADDERS[0].genblk1.FA.sum ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _501_ (.A(\BLOCKS[1].ADDERS[1].genblk1.FA.sum ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _502_ (.A(\BLOCKS[1].ADDERS[2].genblk1.FA.sum ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _503_ (.A(\BLOCKS[1].ADDERS[3].genblk1.FA.sum ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _504_ (.A(\BLOCKS[2].ADDERS[0].genblk1.FA.sum ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _505_ (.A(\BLOCKS[2].ADDERS[1].genblk1.FA.sum ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _506_ (.A(\BLOCKS[2].ADDERS[2].genblk1.FA.sum ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _507_ (.A(\BLOCKS[2].ADDERS[3].genblk1.FA.sum ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _508_ (.A(\BLOCKS[3].ADDERS[0].genblk1.FA.sum ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _509_ (.A(\BLOCKS[3].ADDERS[1].genblk1.FA.sum ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _510_ (.A(\BLOCKS[3].ADDERS[2].genblk1.FA.sum ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _511_ (.A(\BLOCKS[3].ADDERS[3].genblk1.FA.sum ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _512_ (.A(\BLOCKS[4].ADDERS[0].genblk1.FA.sum ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _513_ (.A(\BLOCKS[4].ADDERS[1].genblk1.FA.sum ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _514_ (.A(\BLOCKS[4].ADDERS[2].genblk1.FA.sum ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _515_ (.A(\BLOCKS[4].ADDERS[3].genblk1.FA.sum ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _516_ (.A(\BLOCKS[5].ADDERS[0].genblk1.FA.sum ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _517_ (.A(\BLOCKS[5].ADDERS[1].genblk1.FA.sum ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _518_ (.A(\BLOCKS[5].ADDERS[2].genblk1.FA.sum ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _519_ (.A(\BLOCKS[5].ADDERS[3].genblk1.FA.sum ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _520_ (.A(\BLOCKS[6].ADDERS[0].genblk1.FA.sum ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _521_ (.A(\BLOCKS[6].ADDERS[1].genblk1.FA.sum ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _522_ (.A(\BLOCKS[6].ADDERS[2].genblk1.FA.sum ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _523_ (.A(\BLOCKS[6].ADDERS[3].genblk1.FA.sum ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _524_ (.A(\BLOCKS[7].ADDERS[0].genblk1.FA.sum ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _525_ (.A(\BLOCKS[7].ADDERS[1].genblk1.FA.sum ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _526_ (.A(\BLOCKS[7].ADDERS[2].genblk1.FA.sum ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _527_ (.A(\BLOCKS[7].ADDERS[3].genblk1.FA.sum ),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(Cin),
    .X(net65));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(Cout));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(Overflow));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(Sum[0]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(Sum[10]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(Sum[11]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(Sum[12]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(Sum[13]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(Sum[14]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(Sum[15]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(Sum[16]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(Sum[17]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(Sum[18]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(Sum[19]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(Sum[1]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(Sum[20]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(Sum[21]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(Sum[22]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(Sum[23]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(Sum[24]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(Sum[25]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(Sum[26]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(Sum[27]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(Sum[28]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(Sum[29]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(Sum[2]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(Sum[30]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(Sum[31]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(Sum[3]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(Sum[4]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(Sum[5]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(Sum[6]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(Sum[7]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(Sum[8]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(Sum[9]));
endmodule
