module CarrySelectAdder (Cin,
    Cout,
    Overflow,
    A,
    B,
    Sum);
 input Cin;
 output Cout;
 output Overflow;
 input [31:0] A;
 input [31:0] B;
 output [31:0] Sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__inv_2 _166_ (.A(net55),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _167_ (.A(net23),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_1 _168_ (.A(net33),
    .B(net1),
    .Y(_002_));
 sky130_fd_sc_hd__and3_1 _169_ (.A(net65),
    .B(net33),
    .C(net1),
    .X(_003_));
 sky130_fd_sc_hd__or2_1 _170_ (.A(net33),
    .B(net1),
    .X(_004_));
 sky130_fd_sc_hd__o21ai_1 _171_ (.A1(net33),
    .A2(net1),
    .B1(net65),
    .Y(_005_));
 sky130_fd_sc_hd__and2_1 _172_ (.A(_002_),
    .B(_005_),
    .X(_006_));
 sky130_fd_sc_hd__o22a_1 _173_ (.A1(_004_),
    .A2(net65),
    .B1(_003_),
    .B2(_006_),
    .X(net68));
 sky130_fd_sc_hd__nor2_1 _174_ (.A(net57),
    .B(net25),
    .Y(_007_));
 sky130_fd_sc_hd__or2_1 _175_ (.A(net57),
    .B(net25),
    .X(_008_));
 sky130_fd_sc_hd__and2_1 _176_ (.A(net57),
    .B(net25),
    .X(_009_));
 sky130_fd_sc_hd__nand2_1 _177_ (.A(net57),
    .B(net25),
    .Y(_010_));
 sky130_fd_sc_hd__and2_1 _178_ (.A(net56),
    .B(net24),
    .X(_011_));
 sky130_fd_sc_hd__nand2_1 _179_ (.A(net56),
    .B(net24),
    .Y(_012_));
 sky130_fd_sc_hd__and2_1 _180_ (.A(net54),
    .B(net22),
    .X(_013_));
 sky130_fd_sc_hd__nor2_1 _181_ (.A(net54),
    .B(net22),
    .Y(_014_));
 sky130_fd_sc_hd__nor2_1 _182_ (.A(_013_),
    .B(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__and2_1 _183_ (.A(net53),
    .B(net21),
    .X(_016_));
 sky130_fd_sc_hd__and2_1 _184_ (.A(net52),
    .B(net20),
    .X(_017_));
 sky130_fd_sc_hd__nor2_1 _185_ (.A(net52),
    .B(net20),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_1 _186_ (.A(_017_),
    .B(_018_),
    .Y(_019_));
 sky130_fd_sc_hd__and2_1 _187_ (.A(net51),
    .B(net19),
    .X(_020_));
 sky130_fd_sc_hd__and2_1 _188_ (.A(net50),
    .B(net18),
    .X(_021_));
 sky130_fd_sc_hd__nor2_1 _189_ (.A(net50),
    .B(net18),
    .Y(_022_));
 sky130_fd_sc_hd__nor2_1 _190_ (.A(_021_),
    .B(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__and2_1 _191_ (.A(net49),
    .B(net17),
    .X(_024_));
 sky130_fd_sc_hd__and2_1 _192_ (.A(net48),
    .B(net16),
    .X(_025_));
 sky130_fd_sc_hd__nor2_1 _193_ (.A(net48),
    .B(net16),
    .Y(_026_));
 sky130_fd_sc_hd__nor2_1 _194_ (.A(_025_),
    .B(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__and2_1 _195_ (.A(net47),
    .B(net15),
    .X(_028_));
 sky130_fd_sc_hd__and2_1 _196_ (.A(net46),
    .B(net14),
    .X(_029_));
 sky130_fd_sc_hd__nor2_1 _197_ (.A(net46),
    .B(net14),
    .Y(_030_));
 sky130_fd_sc_hd__nor2_1 _198_ (.A(_029_),
    .B(_030_),
    .Y(_031_));
 sky130_fd_sc_hd__and2_1 _199_ (.A(net45),
    .B(net13),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _200_ (.A(net43),
    .B(net11),
    .X(_033_));
 sky130_fd_sc_hd__nor2_1 _201_ (.A(net43),
    .B(net11),
    .Y(_034_));
 sky130_fd_sc_hd__nor2_1 _202_ (.A(_033_),
    .B(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__and2_1 _203_ (.A(net42),
    .B(net10),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _204_ (.A(net41),
    .B(net9),
    .X(_037_));
 sky130_fd_sc_hd__nor2_1 _205_ (.A(net41),
    .B(net9),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _206_ (.A(_037_),
    .B(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__and2_1 _207_ (.A(net40),
    .B(net8),
    .X(_040_));
 sky130_fd_sc_hd__and2_1 _208_ (.A(net39),
    .B(net7),
    .X(_041_));
 sky130_fd_sc_hd__nor2_1 _209_ (.A(net39),
    .B(net7),
    .Y(_042_));
 sky130_fd_sc_hd__nor2_1 _210_ (.A(_041_),
    .B(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__and2_1 _211_ (.A(net38),
    .B(net6),
    .X(_044_));
 sky130_fd_sc_hd__and2_1 _212_ (.A(net37),
    .B(net5),
    .X(_045_));
 sky130_fd_sc_hd__nor2_1 _213_ (.A(net37),
    .B(net5),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_1 _214_ (.A(_045_),
    .B(_046_),
    .Y(_047_));
 sky130_fd_sc_hd__and2_1 _215_ (.A(net36),
    .B(net4),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _216_ (.A(net35),
    .B(net3),
    .X(_049_));
 sky130_fd_sc_hd__nor2_1 _217_ (.A(net35),
    .B(net3),
    .Y(_050_));
 sky130_fd_sc_hd__nor2_1 _218_ (.A(_049_),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__and2_1 _219_ (.A(net34),
    .B(net2),
    .X(_052_));
 sky130_fd_sc_hd__and2_1 _220_ (.A(net64),
    .B(net32),
    .X(_053_));
 sky130_fd_sc_hd__nor2_1 _221_ (.A(net64),
    .B(net32),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _222_ (.A(_053_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__and2_1 _223_ (.A(net63),
    .B(net31),
    .X(_056_));
 sky130_fd_sc_hd__and2_1 _224_ (.A(net62),
    .B(net30),
    .X(_057_));
 sky130_fd_sc_hd__nor2_1 _225_ (.A(net62),
    .B(net30),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _226_ (.A(_057_),
    .B(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__and2_1 _227_ (.A(net61),
    .B(net29),
    .X(_060_));
 sky130_fd_sc_hd__and2_1 _228_ (.A(net60),
    .B(net28),
    .X(_061_));
 sky130_fd_sc_hd__nor2_1 _229_ (.A(net60),
    .B(net28),
    .Y(_062_));
 sky130_fd_sc_hd__nor2_1 _230_ (.A(_061_),
    .B(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__and2_1 _231_ (.A(net59),
    .B(net27),
    .X(_064_));
 sky130_fd_sc_hd__and2_1 _232_ (.A(net58),
    .B(net26),
    .X(_065_));
 sky130_fd_sc_hd__nor2_1 _233_ (.A(net58),
    .B(net26),
    .Y(_066_));
 sky130_fd_sc_hd__nor2_1 _234_ (.A(_065_),
    .B(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__nor2_1 _235_ (.A(_000_),
    .B(_001_),
    .Y(_068_));
 sky130_fd_sc_hd__nand2_1 _236_ (.A(net55),
    .B(net23),
    .Y(_069_));
 sky130_fd_sc_hd__or2_1 _237_ (.A(net55),
    .B(net23),
    .X(_070_));
 sky130_fd_sc_hd__or2_1 _238_ (.A(net44),
    .B(net12),
    .X(_071_));
 sky130_fd_sc_hd__nand2_1 _239_ (.A(net44),
    .B(net12),
    .Y(_072_));
 sky130_fd_sc_hd__nand3_1 _240_ (.A(_002_),
    .B(_005_),
    .C(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__o2111ai_1 _241_ (.A1(net44),
    .A2(net12),
    .B1(_069_),
    .C1(_070_),
    .D1(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__a31oi_2 _242_ (.A1(_070_),
    .A2(_071_),
    .A3(_073_),
    .B1(_068_),
    .Y(_075_));
 sky130_fd_sc_hd__o21ai_1 _243_ (.A1(_000_),
    .A2(_001_),
    .B1(_074_),
    .Y(_076_));
 sky130_fd_sc_hd__a21oi_1 _244_ (.A1(_076_),
    .A2(_067_),
    .B1(_065_),
    .Y(_077_));
 sky130_fd_sc_hd__o21bai_1 _245_ (.A1(_066_),
    .A2(_075_),
    .B1_N(_065_),
    .Y(_078_));
 sky130_fd_sc_hd__or2_1 _246_ (.A(net59),
    .B(net27),
    .X(_079_));
 sky130_fd_sc_hd__nand2b_1 _247_ (.A_N(_064_),
    .B(_079_),
    .Y(_080_));
 sky130_fd_sc_hd__a21oi_1 _248_ (.A1(_078_),
    .A2(_079_),
    .B1(_064_),
    .Y(_081_));
 sky130_fd_sc_hd__o21bai_1 _249_ (.A1(_080_),
    .A2(_077_),
    .B1_N(_064_),
    .Y(_082_));
 sky130_fd_sc_hd__a21oi_1 _250_ (.A1(_082_),
    .A2(_063_),
    .B1(_061_),
    .Y(_083_));
 sky130_fd_sc_hd__o21bai_1 _251_ (.A1(_062_),
    .A2(_081_),
    .B1_N(_061_),
    .Y(_084_));
 sky130_fd_sc_hd__or2_1 _252_ (.A(net61),
    .B(net29),
    .X(_085_));
 sky130_fd_sc_hd__nand2b_1 _253_ (.A_N(_060_),
    .B(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__a21oi_1 _254_ (.A1(_084_),
    .A2(_085_),
    .B1(_060_),
    .Y(_087_));
 sky130_fd_sc_hd__o21bai_1 _255_ (.A1(_086_),
    .A2(_083_),
    .B1_N(_060_),
    .Y(_088_));
 sky130_fd_sc_hd__a21oi_1 _256_ (.A1(_088_),
    .A2(_059_),
    .B1(_057_),
    .Y(_089_));
 sky130_fd_sc_hd__o21bai_1 _257_ (.A1(_058_),
    .A2(_087_),
    .B1_N(_057_),
    .Y(_090_));
 sky130_fd_sc_hd__or2_1 _258_ (.A(net63),
    .B(net31),
    .X(_091_));
 sky130_fd_sc_hd__nand2b_1 _259_ (.A_N(_056_),
    .B(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__a21oi_1 _260_ (.A1(_090_),
    .A2(_091_),
    .B1(_056_),
    .Y(_093_));
 sky130_fd_sc_hd__o21bai_1 _261_ (.A1(_092_),
    .A2(_089_),
    .B1_N(_056_),
    .Y(_094_));
 sky130_fd_sc_hd__a21oi_1 _262_ (.A1(_094_),
    .A2(_055_),
    .B1(_053_),
    .Y(_095_));
 sky130_fd_sc_hd__o21bai_2 _263_ (.A1(_054_),
    .A2(_093_),
    .B1_N(_053_),
    .Y(_096_));
 sky130_fd_sc_hd__or2_1 _264_ (.A(net34),
    .B(net2),
    .X(_097_));
 sky130_fd_sc_hd__nand2b_1 _265_ (.A_N(_052_),
    .B(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__a21oi_1 _266_ (.A1(_096_),
    .A2(_097_),
    .B1(_052_),
    .Y(_099_));
 sky130_fd_sc_hd__o21bai_1 _267_ (.A1(_098_),
    .A2(_095_),
    .B1_N(_052_),
    .Y(_100_));
 sky130_fd_sc_hd__a21oi_1 _268_ (.A1(_100_),
    .A2(_051_),
    .B1(_049_),
    .Y(_101_));
 sky130_fd_sc_hd__o21bai_2 _269_ (.A1(_050_),
    .A2(_099_),
    .B1_N(_049_),
    .Y(_102_));
 sky130_fd_sc_hd__or2_1 _270_ (.A(net36),
    .B(net4),
    .X(_103_));
 sky130_fd_sc_hd__nand2b_1 _271_ (.A_N(_048_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__a21oi_1 _272_ (.A1(_102_),
    .A2(_103_),
    .B1(_048_),
    .Y(_105_));
 sky130_fd_sc_hd__o21bai_1 _273_ (.A1(_104_),
    .A2(_101_),
    .B1_N(_048_),
    .Y(_106_));
 sky130_fd_sc_hd__a21oi_1 _274_ (.A1(_106_),
    .A2(_047_),
    .B1(_045_),
    .Y(_107_));
 sky130_fd_sc_hd__o21bai_2 _275_ (.A1(_046_),
    .A2(_105_),
    .B1_N(_045_),
    .Y(_108_));
 sky130_fd_sc_hd__or2_1 _276_ (.A(net38),
    .B(net6),
    .X(_109_));
 sky130_fd_sc_hd__nand2b_1 _277_ (.A_N(_044_),
    .B(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__a21oi_2 _278_ (.A1(_108_),
    .A2(_109_),
    .B1(_044_),
    .Y(_111_));
 sky130_fd_sc_hd__o21bai_1 _279_ (.A1(_110_),
    .A2(_107_),
    .B1_N(_044_),
    .Y(_112_));
 sky130_fd_sc_hd__a21oi_1 _280_ (.A1(_112_),
    .A2(_043_),
    .B1(_041_),
    .Y(_113_));
 sky130_fd_sc_hd__o21bai_4 _281_ (.A1(_042_),
    .A2(_111_),
    .B1_N(_041_),
    .Y(_114_));
 sky130_fd_sc_hd__or2_1 _282_ (.A(net40),
    .B(net8),
    .X(_115_));
 sky130_fd_sc_hd__nand2b_1 _283_ (.A_N(_040_),
    .B(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__a21oi_2 _284_ (.A1(_114_),
    .A2(_115_),
    .B1(_040_),
    .Y(_117_));
 sky130_fd_sc_hd__o21bai_1 _285_ (.A1(_116_),
    .A2(_113_),
    .B1_N(_040_),
    .Y(_118_));
 sky130_fd_sc_hd__a21oi_1 _286_ (.A1(_118_),
    .A2(_039_),
    .B1(_037_),
    .Y(_119_));
 sky130_fd_sc_hd__o21bai_2 _287_ (.A1(_038_),
    .A2(_117_),
    .B1_N(_037_),
    .Y(_120_));
 sky130_fd_sc_hd__or2_1 _288_ (.A(net42),
    .B(net10),
    .X(_121_));
 sky130_fd_sc_hd__nand2b_1 _289_ (.A_N(_036_),
    .B(_121_),
    .Y(_122_));
 sky130_fd_sc_hd__a21oi_1 _290_ (.A1(_120_),
    .A2(_121_),
    .B1(_036_),
    .Y(_123_));
 sky130_fd_sc_hd__o21bai_1 _291_ (.A1(_122_),
    .A2(_119_),
    .B1_N(_036_),
    .Y(_124_));
 sky130_fd_sc_hd__a21oi_1 _292_ (.A1(_124_),
    .A2(_035_),
    .B1(_033_),
    .Y(_125_));
 sky130_fd_sc_hd__o21bai_1 _293_ (.A1(_034_),
    .A2(_123_),
    .B1_N(_033_),
    .Y(_126_));
 sky130_fd_sc_hd__or2_1 _294_ (.A(net45),
    .B(net13),
    .X(_127_));
 sky130_fd_sc_hd__nand2b_1 _295_ (.A_N(_032_),
    .B(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__a21oi_1 _296_ (.A1(_126_),
    .A2(_127_),
    .B1(_032_),
    .Y(_129_));
 sky130_fd_sc_hd__o21bai_1 _297_ (.A1(_128_),
    .A2(_125_),
    .B1_N(_032_),
    .Y(_130_));
 sky130_fd_sc_hd__a21oi_1 _298_ (.A1(_130_),
    .A2(_031_),
    .B1(_029_),
    .Y(_131_));
 sky130_fd_sc_hd__o21bai_1 _299_ (.A1(_030_),
    .A2(_129_),
    .B1_N(_029_),
    .Y(_132_));
 sky130_fd_sc_hd__or2_1 _300_ (.A(net47),
    .B(net15),
    .X(_133_));
 sky130_fd_sc_hd__nand2b_1 _301_ (.A_N(_028_),
    .B(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__a21oi_1 _302_ (.A1(_132_),
    .A2(_133_),
    .B1(_028_),
    .Y(_135_));
 sky130_fd_sc_hd__o21bai_1 _303_ (.A1(_134_),
    .A2(_131_),
    .B1_N(_028_),
    .Y(_136_));
 sky130_fd_sc_hd__a21oi_1 _304_ (.A1(_136_),
    .A2(_027_),
    .B1(_025_),
    .Y(_137_));
 sky130_fd_sc_hd__o21bai_1 _305_ (.A1(_026_),
    .A2(_135_),
    .B1_N(_025_),
    .Y(_138_));
 sky130_fd_sc_hd__or2_1 _306_ (.A(net49),
    .B(net17),
    .X(_139_));
 sky130_fd_sc_hd__nand2b_1 _307_ (.A_N(_024_),
    .B(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__a21oi_1 _308_ (.A1(_138_),
    .A2(_139_),
    .B1(_024_),
    .Y(_141_));
 sky130_fd_sc_hd__o21bai_1 _309_ (.A1(_140_),
    .A2(_137_),
    .B1_N(_024_),
    .Y(_142_));
 sky130_fd_sc_hd__a21oi_1 _310_ (.A1(_142_),
    .A2(_023_),
    .B1(_021_),
    .Y(_143_));
 sky130_fd_sc_hd__o21bai_1 _311_ (.A1(_022_),
    .A2(_141_),
    .B1_N(_021_),
    .Y(_144_));
 sky130_fd_sc_hd__or2_1 _312_ (.A(net51),
    .B(net19),
    .X(_145_));
 sky130_fd_sc_hd__nand2b_1 _313_ (.A_N(_020_),
    .B(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__a21oi_1 _314_ (.A1(_144_),
    .A2(_145_),
    .B1(_020_),
    .Y(_147_));
 sky130_fd_sc_hd__o21bai_1 _315_ (.A1(_146_),
    .A2(_143_),
    .B1_N(_020_),
    .Y(_148_));
 sky130_fd_sc_hd__a21oi_1 _316_ (.A1(_148_),
    .A2(_019_),
    .B1(_017_),
    .Y(_149_));
 sky130_fd_sc_hd__o21bai_2 _317_ (.A1(_018_),
    .A2(_147_),
    .B1_N(_017_),
    .Y(_150_));
 sky130_fd_sc_hd__or2_1 _318_ (.A(net53),
    .B(net21),
    .X(_151_));
 sky130_fd_sc_hd__nand2b_1 _319_ (.A_N(_016_),
    .B(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__a21oi_2 _320_ (.A1(_150_),
    .A2(_151_),
    .B1(_016_),
    .Y(_153_));
 sky130_fd_sc_hd__o21bai_1 _321_ (.A1(_152_),
    .A2(_149_),
    .B1_N(_016_),
    .Y(_154_));
 sky130_fd_sc_hd__a21oi_1 _322_ (.A1(_154_),
    .A2(_015_),
    .B1(_013_),
    .Y(_155_));
 sky130_fd_sc_hd__o21bai_1 _323_ (.A1(_014_),
    .A2(_153_),
    .B1_N(_013_),
    .Y(_156_));
 sky130_fd_sc_hd__or2_1 _324_ (.A(net56),
    .B(net24),
    .X(_157_));
 sky130_fd_sc_hd__nand2_1 _325_ (.A(_012_),
    .B(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__a21oi_1 _326_ (.A1(_156_),
    .A2(_157_),
    .B1(_011_),
    .Y(_159_));
 sky130_fd_sc_hd__o21bai_1 _327_ (.A1(_158_),
    .A2(_155_),
    .B1_N(_011_),
    .Y(_160_));
 sky130_fd_sc_hd__o21ai_1 _328_ (.A1(_007_),
    .A2(_009_),
    .B1(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__o2111ai_1 _329_ (.A1(_158_),
    .A2(_155_),
    .B1(_010_),
    .C1(_008_),
    .D1(_012_),
    .Y(_162_));
 sky130_fd_sc_hd__nand2_1 _330_ (.A(_161_),
    .B(_162_),
    .Y(net92));
 sky130_fd_sc_hd__o211ai_1 _331_ (.A1(_158_),
    .A2(_155_),
    .B1(_012_),
    .C1(_010_),
    .Y(_163_));
 sky130_fd_sc_hd__o21a_1 _332_ (.A1(_007_),
    .A2(_159_),
    .B1(_163_),
    .X(net67));
 sky130_fd_sc_hd__nand2_1 _333_ (.A(_071_),
    .B(_072_),
    .Y(_164_));
 sky130_fd_sc_hd__xor2_2 _334_ (.A(_006_),
    .B(_164_),
    .X(net79));
 sky130_fd_sc_hd__a22o_1 _335_ (.A1(_069_),
    .A2(_070_),
    .B1(_071_),
    .B2(_073_),
    .X(_165_));
 sky130_fd_sc_hd__and2_1 _336_ (.A(_074_),
    .B(_165_),
    .X(net90));
 sky130_fd_sc_hd__xnor2_1 _337_ (.A(_067_),
    .B(_075_),
    .Y(net93));
 sky130_fd_sc_hd__xnor2_1 _338_ (.A(_078_),
    .B(_080_),
    .Y(net94));
 sky130_fd_sc_hd__xnor2_1 _339_ (.A(_063_),
    .B(_081_),
    .Y(net95));
 sky130_fd_sc_hd__xnor2_1 _340_ (.A(_084_),
    .B(_086_),
    .Y(net96));
 sky130_fd_sc_hd__xnor2_1 _341_ (.A(_059_),
    .B(_087_),
    .Y(net97));
 sky130_fd_sc_hd__xnor2_1 _342_ (.A(_090_),
    .B(_092_),
    .Y(net98));
 sky130_fd_sc_hd__xnor2_1 _343_ (.A(_055_),
    .B(_093_),
    .Y(net99));
 sky130_fd_sc_hd__xnor2_2 _344_ (.A(_096_),
    .B(_098_),
    .Y(net69));
 sky130_fd_sc_hd__xnor2_1 _345_ (.A(_051_),
    .B(_099_),
    .Y(net70));
 sky130_fd_sc_hd__xnor2_1 _346_ (.A(_102_),
    .B(_104_),
    .Y(net71));
 sky130_fd_sc_hd__xnor2_1 _347_ (.A(_047_),
    .B(_105_),
    .Y(net72));
 sky130_fd_sc_hd__xnor2_1 _348_ (.A(_108_),
    .B(_110_),
    .Y(net73));
 sky130_fd_sc_hd__xnor2_1 _349_ (.A(_043_),
    .B(_111_),
    .Y(net74));
 sky130_fd_sc_hd__xnor2_2 _350_ (.A(_114_),
    .B(_116_),
    .Y(net75));
 sky130_fd_sc_hd__xnor2_2 _351_ (.A(_039_),
    .B(_117_),
    .Y(net76));
 sky130_fd_sc_hd__xnor2_2 _352_ (.A(_120_),
    .B(_122_),
    .Y(net77));
 sky130_fd_sc_hd__xnor2_1 _353_ (.A(_035_),
    .B(_123_),
    .Y(net78));
 sky130_fd_sc_hd__xnor2_1 _354_ (.A(_126_),
    .B(_128_),
    .Y(net80));
 sky130_fd_sc_hd__xnor2_1 _355_ (.A(_031_),
    .B(_129_),
    .Y(net81));
 sky130_fd_sc_hd__xnor2_1 _356_ (.A(_132_),
    .B(_134_),
    .Y(net82));
 sky130_fd_sc_hd__xnor2_1 _357_ (.A(_027_),
    .B(_135_),
    .Y(net83));
 sky130_fd_sc_hd__xnor2_1 _358_ (.A(_138_),
    .B(_140_),
    .Y(net84));
 sky130_fd_sc_hd__xnor2_1 _359_ (.A(_023_),
    .B(_141_),
    .Y(net85));
 sky130_fd_sc_hd__xnor2_1 _360_ (.A(_144_),
    .B(_146_),
    .Y(net86));
 sky130_fd_sc_hd__xnor2_1 _361_ (.A(_019_),
    .B(_147_),
    .Y(net87));
 sky130_fd_sc_hd__xnor2_1 _362_ (.A(_150_),
    .B(_152_),
    .Y(net88));
 sky130_fd_sc_hd__xnor2_2 _363_ (.A(_015_),
    .B(_153_),
    .Y(net89));
 sky130_fd_sc_hd__xnor2_1 _364_ (.A(_156_),
    .B(_158_),
    .Y(net91));
 sky130_fd_sc_hd__a21oi_1 _365_ (.A1(_159_),
    .A2(_010_),
    .B1(_007_),
    .Y(net66));
 sky130_fd_sc_hd__buf_1 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(Cin),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 output66 (.A(net66),
    .X(Cout));
 sky130_fd_sc_hd__clkbuf_16 output67 (.A(net67),
    .X(Overflow));
 sky130_fd_sc_hd__clkbuf_16 output68 (.A(net68),
    .X(Sum[0]));
 sky130_fd_sc_hd__clkbuf_16 output69 (.A(net69),
    .X(Sum[10]));
 sky130_fd_sc_hd__clkbuf_16 output70 (.A(net70),
    .X(Sum[11]));
 sky130_fd_sc_hd__clkbuf_16 output71 (.A(net71),
    .X(Sum[12]));
 sky130_fd_sc_hd__clkbuf_16 output72 (.A(net72),
    .X(Sum[13]));
 sky130_fd_sc_hd__clkbuf_16 output73 (.A(net73),
    .X(Sum[14]));
 sky130_fd_sc_hd__clkbuf_16 output74 (.A(net74),
    .X(Sum[15]));
 sky130_fd_sc_hd__clkbuf_16 output75 (.A(net75),
    .X(Sum[16]));
 sky130_fd_sc_hd__clkbuf_16 output76 (.A(net76),
    .X(Sum[17]));
 sky130_fd_sc_hd__clkbuf_16 output77 (.A(net77),
    .X(Sum[18]));
 sky130_fd_sc_hd__clkbuf_16 output78 (.A(net78),
    .X(Sum[19]));
 sky130_fd_sc_hd__clkbuf_16 output79 (.A(net79),
    .X(Sum[1]));
 sky130_fd_sc_hd__clkbuf_16 output80 (.A(net80),
    .X(Sum[20]));
 sky130_fd_sc_hd__clkbuf_16 output81 (.A(net81),
    .X(Sum[21]));
 sky130_fd_sc_hd__clkbuf_16 output82 (.A(net82),
    .X(Sum[22]));
 sky130_fd_sc_hd__clkbuf_16 output83 (.A(net83),
    .X(Sum[23]));
 sky130_fd_sc_hd__clkbuf_16 output84 (.A(net84),
    .X(Sum[24]));
 sky130_fd_sc_hd__clkbuf_16 output85 (.A(net85),
    .X(Sum[25]));
 sky130_fd_sc_hd__clkbuf_16 output86 (.A(net86),
    .X(Sum[26]));
 sky130_fd_sc_hd__clkbuf_16 output87 (.A(net87),
    .X(Sum[27]));
 sky130_fd_sc_hd__clkbuf_16 output88 (.A(net88),
    .X(Sum[28]));
 sky130_fd_sc_hd__clkbuf_16 output89 (.A(net89),
    .X(Sum[29]));
 sky130_fd_sc_hd__clkbuf_16 output90 (.A(net90),
    .X(Sum[2]));
 sky130_fd_sc_hd__clkbuf_16 output91 (.A(net91),
    .X(Sum[30]));
 sky130_fd_sc_hd__clkbuf_16 output92 (.A(net92),
    .X(Sum[31]));
 sky130_fd_sc_hd__clkbuf_16 output93 (.A(net93),
    .X(Sum[3]));
 sky130_fd_sc_hd__clkbuf_16 output94 (.A(net94),
    .X(Sum[4]));
 sky130_fd_sc_hd__clkbuf_16 output95 (.A(net95),
    .X(Sum[5]));
 sky130_fd_sc_hd__clkbuf_16 output96 (.A(net96),
    .X(Sum[6]));
 sky130_fd_sc_hd__clkbuf_16 output97 (.A(net97),
    .X(Sum[7]));
 sky130_fd_sc_hd__clkbuf_16 output98 (.A(net98),
    .X(Sum[8]));
 sky130_fd_sc_hd__clkbuf_16 output99 (.A(net99),
    .X(Sum[9]));
endmodule
