module ripple_carry_adder (overflow,
    a,
    b,
    sum);
 output overflow;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire \FA0.p1 ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire \ripple[10].FA.sum ;
 wire \ripple[11].FA.sum ;
 wire \ripple[12].FA.sum ;
 wire \ripple[13].FA.sum ;
 wire \ripple[14].FA.sum ;
 wire \ripple[15].FA.sum ;
 wire \ripple[16].FA.sum ;
 wire \ripple[17].FA.sum ;
 wire \ripple[18].FA.sum ;
 wire \ripple[19].FA.sum ;
 wire \ripple[1].FA.sum ;
 wire \ripple[20].FA.sum ;
 wire \ripple[21].FA.sum ;
 wire \ripple[22].FA.sum ;
 wire \ripple[23].FA.sum ;
 wire \ripple[24].FA.sum ;
 wire \ripple[25].FA.sum ;
 wire \ripple[26].FA.sum ;
 wire \ripple[27].FA.sum ;
 wire \ripple[28].FA.sum ;
 wire \ripple[29].FA.sum ;
 wire \ripple[2].FA.sum ;
 wire \ripple[30].FA.sum ;
 wire \ripple[31].FA.sum ;
 wire \ripple[3].FA.sum ;
 wire \ripple[4].FA.sum ;
 wire \ripple[5].FA.sum ;
 wire \ripple[6].FA.sum ;
 wire \ripple[7].FA.sum ;
 wire \ripple[8].FA.sum ;
 wire \ripple[9].FA.sum ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;

 sky130_fd_sc_hd__nor2_1 _133_ (.A(net57),
    .B(net25),
    .Y(_131_));
 sky130_fd_sc_hd__or2_1 _134_ (.A(net57),
    .B(net25),
    .X(_132_));
 sky130_fd_sc_hd__and2_1 _135_ (.A(net57),
    .B(net25),
    .X(_000_));
 sky130_fd_sc_hd__nand2_1 _136_ (.A(net57),
    .B(net25),
    .Y(_001_));
 sky130_fd_sc_hd__and2_1 _137_ (.A(net56),
    .B(net24),
    .X(_002_));
 sky130_fd_sc_hd__nand2_1 _138_ (.A(net56),
    .B(net24),
    .Y(_003_));
 sky130_fd_sc_hd__and2_1 _139_ (.A(net54),
    .B(net22),
    .X(_004_));
 sky130_fd_sc_hd__nor2_1 _140_ (.A(net54),
    .B(net22),
    .Y(_005_));
 sky130_fd_sc_hd__nor2_1 _141_ (.A(_004_),
    .B(_005_),
    .Y(_006_));
 sky130_fd_sc_hd__and2_1 _142_ (.A(net53),
    .B(net21),
    .X(_007_));
 sky130_fd_sc_hd__and2_1 _143_ (.A(net52),
    .B(net20),
    .X(_008_));
 sky130_fd_sc_hd__nor2_1 _144_ (.A(net52),
    .B(net20),
    .Y(_009_));
 sky130_fd_sc_hd__nor2_1 _145_ (.A(_008_),
    .B(_009_),
    .Y(_010_));
 sky130_fd_sc_hd__and2_1 _146_ (.A(net51),
    .B(net19),
    .X(_011_));
 sky130_fd_sc_hd__and2_1 _147_ (.A(net50),
    .B(net18),
    .X(_012_));
 sky130_fd_sc_hd__nor2_1 _148_ (.A(net50),
    .B(net18),
    .Y(_013_));
 sky130_fd_sc_hd__nor2_1 _149_ (.A(_012_),
    .B(_013_),
    .Y(_014_));
 sky130_fd_sc_hd__and2_1 _150_ (.A(net49),
    .B(net17),
    .X(_015_));
 sky130_fd_sc_hd__and2_1 _151_ (.A(net48),
    .B(net16),
    .X(_016_));
 sky130_fd_sc_hd__nor2_1 _152_ (.A(net48),
    .B(net16),
    .Y(_017_));
 sky130_fd_sc_hd__nor2_1 _153_ (.A(_016_),
    .B(_017_),
    .Y(_018_));
 sky130_fd_sc_hd__and2_1 _154_ (.A(net47),
    .B(net15),
    .X(_019_));
 sky130_fd_sc_hd__and2_1 _155_ (.A(net46),
    .B(net14),
    .X(_020_));
 sky130_fd_sc_hd__nor2_1 _156_ (.A(net46),
    .B(net14),
    .Y(_021_));
 sky130_fd_sc_hd__nor2_1 _157_ (.A(_020_),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__and2_1 _158_ (.A(net45),
    .B(net13),
    .X(_023_));
 sky130_fd_sc_hd__and2_1 _159_ (.A(net43),
    .B(net11),
    .X(_024_));
 sky130_fd_sc_hd__nor2_1 _160_ (.A(net43),
    .B(net11),
    .Y(_025_));
 sky130_fd_sc_hd__nor2_1 _161_ (.A(_024_),
    .B(_025_),
    .Y(_026_));
 sky130_fd_sc_hd__and2_1 _162_ (.A(net42),
    .B(net10),
    .X(_027_));
 sky130_fd_sc_hd__and2_1 _163_ (.A(net41),
    .B(net9),
    .X(_028_));
 sky130_fd_sc_hd__nor2_1 _164_ (.A(net41),
    .B(net9),
    .Y(_029_));
 sky130_fd_sc_hd__nor2_1 _165_ (.A(_028_),
    .B(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__and2_1 _166_ (.A(net40),
    .B(net8),
    .X(_031_));
 sky130_fd_sc_hd__and2_1 _167_ (.A(net39),
    .B(net7),
    .X(_032_));
 sky130_fd_sc_hd__nor2_1 _168_ (.A(net39),
    .B(net7),
    .Y(_033_));
 sky130_fd_sc_hd__nor2_1 _169_ (.A(_032_),
    .B(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__and2_1 _170_ (.A(net38),
    .B(net6),
    .X(_035_));
 sky130_fd_sc_hd__and2_1 _171_ (.A(net37),
    .B(net5),
    .X(_036_));
 sky130_fd_sc_hd__nor2_1 _172_ (.A(net37),
    .B(net5),
    .Y(_037_));
 sky130_fd_sc_hd__nor2_1 _173_ (.A(_036_),
    .B(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__and2_1 _174_ (.A(net36),
    .B(net4),
    .X(_039_));
 sky130_fd_sc_hd__and2_1 _175_ (.A(net35),
    .B(net3),
    .X(_040_));
 sky130_fd_sc_hd__nor2_1 _176_ (.A(net35),
    .B(net3),
    .Y(_041_));
 sky130_fd_sc_hd__nor2_1 _177_ (.A(_040_),
    .B(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__and2_1 _178_ (.A(net34),
    .B(net2),
    .X(_043_));
 sky130_fd_sc_hd__and2_1 _179_ (.A(net64),
    .B(net32),
    .X(_044_));
 sky130_fd_sc_hd__nor2_1 _180_ (.A(net64),
    .B(net32),
    .Y(_045_));
 sky130_fd_sc_hd__nor2_1 _181_ (.A(_044_),
    .B(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__and2_1 _182_ (.A(net63),
    .B(net31),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _183_ (.A(net62),
    .B(net30),
    .X(_048_));
 sky130_fd_sc_hd__nor2_1 _184_ (.A(net62),
    .B(net30),
    .Y(_049_));
 sky130_fd_sc_hd__nor2_1 _185_ (.A(_048_),
    .B(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__and2_1 _186_ (.A(net61),
    .B(net29),
    .X(_051_));
 sky130_fd_sc_hd__and2_1 _187_ (.A(net60),
    .B(net28),
    .X(_052_));
 sky130_fd_sc_hd__nor2_1 _188_ (.A(net60),
    .B(net28),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_1 _189_ (.A(_052_),
    .B(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__and2_1 _190_ (.A(net59),
    .B(net27),
    .X(_055_));
 sky130_fd_sc_hd__and2_1 _191_ (.A(net58),
    .B(net26),
    .X(_056_));
 sky130_fd_sc_hd__nand2_1 _192_ (.A(net58),
    .B(net26),
    .Y(_057_));
 sky130_fd_sc_hd__or2_1 _193_ (.A(net58),
    .B(net26),
    .X(_058_));
 sky130_fd_sc_hd__or2_1 _194_ (.A(net55),
    .B(net23),
    .X(_059_));
 sky130_fd_sc_hd__nand2_1 _195_ (.A(net55),
    .B(net23),
    .Y(_060_));
 sky130_fd_sc_hd__or2_1 _196_ (.A(net44),
    .B(net12),
    .X(_061_));
 sky130_fd_sc_hd__nand2_1 _197_ (.A(net44),
    .B(net12),
    .Y(_062_));
 sky130_fd_sc_hd__o211ai_1 _198_ (.A1(net44),
    .A2(net12),
    .B1(net33),
    .C1(net1),
    .Y(_063_));
 sky130_fd_sc_hd__and2_1 _199_ (.A(_062_),
    .B(_063_),
    .X(_064_));
 sky130_fd_sc_hd__nand3_1 _200_ (.A(_060_),
    .B(_062_),
    .C(_063_),
    .Y(_065_));
 sky130_fd_sc_hd__o2111ai_1 _201_ (.A1(net55),
    .A2(net23),
    .B1(_057_),
    .C1(_058_),
    .D1(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__a31oi_2 _202_ (.A1(_058_),
    .A2(_059_),
    .A3(_065_),
    .B1(_056_),
    .Y(_067_));
 sky130_fd_sc_hd__nor2_1 _203_ (.A(net59),
    .B(net27),
    .Y(_068_));
 sky130_fd_sc_hd__or2_1 _204_ (.A(_055_),
    .B(_068_),
    .X(_069_));
 sky130_fd_sc_hd__o21bai_1 _205_ (.A1(_069_),
    .A2(_067_),
    .B1_N(_055_),
    .Y(_070_));
 sky130_fd_sc_hd__a21oi_1 _206_ (.A1(_070_),
    .A2(_054_),
    .B1(_052_),
    .Y(_071_));
 sky130_fd_sc_hd__nor2_1 _207_ (.A(net61),
    .B(net29),
    .Y(_072_));
 sky130_fd_sc_hd__or2_1 _208_ (.A(_051_),
    .B(_072_),
    .X(_073_));
 sky130_fd_sc_hd__o21bai_1 _209_ (.A1(_073_),
    .A2(_071_),
    .B1_N(_051_),
    .Y(_074_));
 sky130_fd_sc_hd__a21oi_1 _210_ (.A1(_074_),
    .A2(_050_),
    .B1(_048_),
    .Y(_075_));
 sky130_fd_sc_hd__nor2_1 _211_ (.A(net63),
    .B(net31),
    .Y(_076_));
 sky130_fd_sc_hd__or2_1 _212_ (.A(_047_),
    .B(_076_),
    .X(_077_));
 sky130_fd_sc_hd__o21bai_1 _213_ (.A1(_077_),
    .A2(_075_),
    .B1_N(_047_),
    .Y(_078_));
 sky130_fd_sc_hd__a21oi_1 _214_ (.A1(_078_),
    .A2(_046_),
    .B1(_044_),
    .Y(_079_));
 sky130_fd_sc_hd__nor2_1 _215_ (.A(net34),
    .B(net2),
    .Y(_080_));
 sky130_fd_sc_hd__or2_1 _216_ (.A(_043_),
    .B(_080_),
    .X(_081_));
 sky130_fd_sc_hd__o21bai_1 _217_ (.A1(_081_),
    .A2(_079_),
    .B1_N(_043_),
    .Y(_082_));
 sky130_fd_sc_hd__a21oi_1 _218_ (.A1(_082_),
    .A2(_042_),
    .B1(_040_),
    .Y(_083_));
 sky130_fd_sc_hd__nor2_1 _219_ (.A(net36),
    .B(net4),
    .Y(_084_));
 sky130_fd_sc_hd__or2_1 _220_ (.A(_039_),
    .B(_084_),
    .X(_085_));
 sky130_fd_sc_hd__o21bai_2 _221_ (.A1(_085_),
    .A2(_083_),
    .B1_N(_039_),
    .Y(_086_));
 sky130_fd_sc_hd__a21oi_1 _222_ (.A1(_086_),
    .A2(_038_),
    .B1(_036_),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_1 _223_ (.A(net38),
    .B(net6),
    .Y(_088_));
 sky130_fd_sc_hd__or2_1 _224_ (.A(_035_),
    .B(_088_),
    .X(_089_));
 sky130_fd_sc_hd__o21bai_2 _225_ (.A1(_089_),
    .A2(_087_),
    .B1_N(_035_),
    .Y(_090_));
 sky130_fd_sc_hd__a21oi_1 _226_ (.A1(_090_),
    .A2(_034_),
    .B1(_032_),
    .Y(_091_));
 sky130_fd_sc_hd__nor2_1 _227_ (.A(net40),
    .B(net8),
    .Y(_092_));
 sky130_fd_sc_hd__or2_1 _228_ (.A(_031_),
    .B(_092_),
    .X(_093_));
 sky130_fd_sc_hd__o21bai_2 _229_ (.A1(_093_),
    .A2(_091_),
    .B1_N(_031_),
    .Y(_094_));
 sky130_fd_sc_hd__a21oi_2 _230_ (.A1(_094_),
    .A2(_030_),
    .B1(_028_),
    .Y(_095_));
 sky130_fd_sc_hd__nor2_1 _231_ (.A(net42),
    .B(net10),
    .Y(_096_));
 sky130_fd_sc_hd__or2_1 _232_ (.A(_027_),
    .B(_096_),
    .X(_097_));
 sky130_fd_sc_hd__o21bai_1 _233_ (.A1(_097_),
    .A2(_095_),
    .B1_N(_027_),
    .Y(_098_));
 sky130_fd_sc_hd__a21oi_1 _234_ (.A1(_098_),
    .A2(_026_),
    .B1(_024_),
    .Y(_099_));
 sky130_fd_sc_hd__nor2_1 _235_ (.A(net45),
    .B(net13),
    .Y(_100_));
 sky130_fd_sc_hd__or2_1 _236_ (.A(_023_),
    .B(_100_),
    .X(_101_));
 sky130_fd_sc_hd__o21bai_1 _237_ (.A1(_101_),
    .A2(_099_),
    .B1_N(_023_),
    .Y(_102_));
 sky130_fd_sc_hd__a21oi_1 _238_ (.A1(_102_),
    .A2(_022_),
    .B1(_020_),
    .Y(_103_));
 sky130_fd_sc_hd__nor2_1 _239_ (.A(net47),
    .B(net15),
    .Y(_104_));
 sky130_fd_sc_hd__or2_1 _240_ (.A(_019_),
    .B(_104_),
    .X(_105_));
 sky130_fd_sc_hd__o21bai_1 _241_ (.A1(_105_),
    .A2(_103_),
    .B1_N(_019_),
    .Y(_106_));
 sky130_fd_sc_hd__a21oi_1 _242_ (.A1(_106_),
    .A2(_018_),
    .B1(_016_),
    .Y(_107_));
 sky130_fd_sc_hd__nor2_1 _243_ (.A(net49),
    .B(net17),
    .Y(_108_));
 sky130_fd_sc_hd__or2_1 _244_ (.A(_015_),
    .B(_108_),
    .X(_109_));
 sky130_fd_sc_hd__o21bai_1 _245_ (.A1(_109_),
    .A2(_107_),
    .B1_N(_015_),
    .Y(_110_));
 sky130_fd_sc_hd__a21oi_1 _246_ (.A1(_110_),
    .A2(_014_),
    .B1(_012_),
    .Y(_111_));
 sky130_fd_sc_hd__nor2_1 _247_ (.A(net51),
    .B(net19),
    .Y(_112_));
 sky130_fd_sc_hd__or2_1 _248_ (.A(_011_),
    .B(_112_),
    .X(_113_));
 sky130_fd_sc_hd__o21bai_1 _249_ (.A1(_113_),
    .A2(_111_),
    .B1_N(_011_),
    .Y(_114_));
 sky130_fd_sc_hd__a21oi_1 _250_ (.A1(_114_),
    .A2(_010_),
    .B1(_008_),
    .Y(_115_));
 sky130_fd_sc_hd__nor2_1 _251_ (.A(net53),
    .B(net21),
    .Y(_116_));
 sky130_fd_sc_hd__or2_1 _252_ (.A(_007_),
    .B(_116_),
    .X(_117_));
 sky130_fd_sc_hd__o21bai_1 _253_ (.A1(_117_),
    .A2(_115_),
    .B1_N(_007_),
    .Y(_118_));
 sky130_fd_sc_hd__a21oi_2 _254_ (.A1(_118_),
    .A2(_006_),
    .B1(_004_),
    .Y(_119_));
 sky130_fd_sc_hd__or2_1 _255_ (.A(net56),
    .B(net24),
    .X(_120_));
 sky130_fd_sc_hd__nand2_1 _256_ (.A(_003_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__o21bai_1 _257_ (.A1(_121_),
    .A2(_119_),
    .B1_N(_002_),
    .Y(_122_));
 sky130_fd_sc_hd__o2111ai_1 _258_ (.A1(_121_),
    .A2(_119_),
    .B1(_001_),
    .C1(_132_),
    .D1(_003_),
    .Y(_123_));
 sky130_fd_sc_hd__o21ai_1 _259_ (.A1(_131_),
    .A2(_000_),
    .B1(_122_),
    .Y(_124_));
 sky130_fd_sc_hd__nand2_1 _260_ (.A(_123_),
    .B(_124_),
    .Y(\ripple[31].FA.sum ));
 sky130_fd_sc_hd__nand2_1 _261_ (.A(_122_),
    .B(_131_),
    .Y(_125_));
 sky130_fd_sc_hd__o21ai_1 _262_ (.A1(_001_),
    .A2(_122_),
    .B1(_125_),
    .Y(net65));
 sky130_fd_sc_hd__xor2_1 _263_ (.A(net33),
    .B(net1),
    .X(\FA0.p1 ));
 sky130_fd_sc_hd__a22o_1 _264_ (.A1(net33),
    .A2(net1),
    .B1(_061_),
    .B2(_062_),
    .X(_126_));
 sky130_fd_sc_hd__nand4_1 _265_ (.A(_061_),
    .B(_062_),
    .C(net33),
    .D(net1),
    .Y(_127_));
 sky130_fd_sc_hd__and2_1 _266_ (.A(_126_),
    .B(_127_),
    .X(\ripple[1].FA.sum ));
 sky130_fd_sc_hd__a21oi_1 _267_ (.A1(_059_),
    .A2(_060_),
    .B1(_064_),
    .Y(_128_));
 sky130_fd_sc_hd__and3_1 _268_ (.A(_059_),
    .B(_060_),
    .C(_064_),
    .X(_129_));
 sky130_fd_sc_hd__or2_1 _269_ (.A(_128_),
    .B(_129_),
    .X(\ripple[2].FA.sum ));
 sky130_fd_sc_hd__a22o_1 _270_ (.A1(_057_),
    .A2(_058_),
    .B1(_059_),
    .B2(_065_),
    .X(_130_));
 sky130_fd_sc_hd__and2_1 _271_ (.A(_066_),
    .B(_130_),
    .X(\ripple[3].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _272_ (.A(_067_),
    .B(_069_),
    .X(\ripple[4].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _273_ (.A(_054_),
    .B(_070_),
    .X(\ripple[5].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _274_ (.A(_071_),
    .B(_073_),
    .X(\ripple[6].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _275_ (.A(_050_),
    .B(_074_),
    .X(\ripple[7].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _276_ (.A(_075_),
    .B(_077_),
    .X(\ripple[8].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _277_ (.A(_046_),
    .B(_078_),
    .X(\ripple[9].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _278_ (.A(_079_),
    .B(_081_),
    .X(\ripple[10].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _279_ (.A(_042_),
    .B(_082_),
    .X(\ripple[11].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _280_ (.A(_083_),
    .B(_085_),
    .X(\ripple[12].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _281_ (.A(_038_),
    .B(_086_),
    .X(\ripple[13].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _282_ (.A(_087_),
    .B(_089_),
    .X(\ripple[14].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _283_ (.A(_034_),
    .B(_090_),
    .X(\ripple[15].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _284_ (.A(_091_),
    .B(_093_),
    .X(\ripple[16].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _285_ (.A(_030_),
    .B(_094_),
    .X(\ripple[17].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _286_ (.A(_095_),
    .B(_097_),
    .X(\ripple[18].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _287_ (.A(_026_),
    .B(_098_),
    .X(\ripple[19].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _288_ (.A(_099_),
    .B(_101_),
    .X(\ripple[20].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _289_ (.A(_022_),
    .B(_102_),
    .X(\ripple[21].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _290_ (.A(_103_),
    .B(_105_),
    .X(\ripple[22].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _291_ (.A(_018_),
    .B(_106_),
    .X(\ripple[23].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _292_ (.A(_107_),
    .B(_109_),
    .X(\ripple[24].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _293_ (.A(_014_),
    .B(_110_),
    .X(\ripple[25].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _294_ (.A(_111_),
    .B(_113_),
    .X(\ripple[26].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _295_ (.A(_010_),
    .B(_114_),
    .X(\ripple[27].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _296_ (.A(_115_),
    .B(_117_),
    .X(\ripple[28].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _297_ (.A(_006_),
    .B(_118_),
    .X(\ripple[29].FA.sum ));
 sky130_fd_sc_hd__xor2_1 _298_ (.A(_119_),
    .B(_121_),
    .X(\ripple[30].FA.sum ));
 sky130_fd_sc_hd__clkbuf_1 _299_ (.A(\FA0.p1 ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _300_ (.A(\ripple[1].FA.sum ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _301_ (.A(\ripple[2].FA.sum ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _302_ (.A(\ripple[3].FA.sum ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _303_ (.A(\ripple[4].FA.sum ),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _304_ (.A(\ripple[5].FA.sum ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _305_ (.A(\ripple[6].FA.sum ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _306_ (.A(\ripple[7].FA.sum ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _307_ (.A(\ripple[8].FA.sum ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _308_ (.A(\ripple[9].FA.sum ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _309_ (.A(\ripple[10].FA.sum ),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _310_ (.A(\ripple[11].FA.sum ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _311_ (.A(\ripple[12].FA.sum ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _312_ (.A(\ripple[13].FA.sum ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _313_ (.A(\ripple[14].FA.sum ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _314_ (.A(\ripple[15].FA.sum ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _315_ (.A(\ripple[16].FA.sum ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _316_ (.A(\ripple[17].FA.sum ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _317_ (.A(\ripple[18].FA.sum ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _318_ (.A(\ripple[19].FA.sum ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _319_ (.A(\ripple[20].FA.sum ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _320_ (.A(\ripple[21].FA.sum ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _321_ (.A(\ripple[22].FA.sum ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _322_ (.A(\ripple[23].FA.sum ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _323_ (.A(\ripple[24].FA.sum ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _324_ (.A(\ripple[25].FA.sum ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _325_ (.A(\ripple[26].FA.sum ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _326_ (.A(\ripple[27].FA.sum ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _327_ (.A(\ripple[28].FA.sum ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _328_ (.A(\ripple[29].FA.sum ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _329_ (.A(\ripple[30].FA.sum ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _330_ (.A(\ripple[31].FA.sum ),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 output65 (.A(net65),
    .X(overflow));
 sky130_fd_sc_hd__buf_1 output66 (.A(net66),
    .X(sum[0]));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(sum[10]));
 sky130_fd_sc_hd__buf_1 output68 (.A(net68),
    .X(sum[11]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(sum[12]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(sum[13]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(sum[14]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(sum[15]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(sum[16]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(sum[17]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(sum[18]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(sum[19]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(sum[1]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(sum[20]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(sum[21]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(sum[22]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(sum[23]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(sum[24]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(sum[25]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(sum[26]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(sum[27]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(sum[28]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(sum[29]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(sum[2]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(sum[30]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(sum[31]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(sum[3]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(sum[4]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(sum[5]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(sum[6]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(sum[7]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(sum[8]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(sum[9]));
endmodule
